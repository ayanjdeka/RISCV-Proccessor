module dadda_32x32
import mult_funct3::*;
(
    input clk,
    input rst,
    input mult_funct3_t mult_op,
    input logic compute_sign,
    input logic ld_carry,
    //input logic flip_sign,
    input logic mult_done,
    input logic mult_done_flip,
    input logic flip_rs1,
    input logic flip_rs2,
    input logic [31:0] A,
    input logic  [31:0] B,
    output logic  [63:0] C,
    output logic rs1_msb,
    output logic rs2_msb
);

//logic [31:0] pp[32];
logic [19:0] s0, c0;
logic [161:0] s1, c1;
logic [197:0] s2, c2;
logic [171:0] s3, c3;
logic [149:0] s4, c4;
logic [109:0] s5, c5;
logic [57:0]  s6, c6;
logic [59:0]  s7, c7;
logic [61:0] c8;

logic [31:0] A_reg, B_reg;
logic [63:0] C_reg;
logic [63:0] O;
logic carry_31;

assign rs1_msb = A[31];
assign rs2_msb = B[31];

always_ff @(posedge clk) begin: calculate_inputs
    if(rst) begin
        A_reg <= '0;
        B_reg <= '0;
    end
    else if(compute_sign) begin
        if(flip_rs1 && flip_rs2) begin
            A_reg <= ~A + 1;
            B_reg <= ~B + 1;
        end
        else if(flip_rs1) begin
            A_reg <= ~A + 1;
            B_reg <= B;
        end
        else if(flip_rs2) begin
            A_reg <= A;
            B_reg <= ~B + 1;
        end
        else begin
            A_reg <= A;
            B_reg <= B;
        end 
    end
end

// always_ff @ (posedge clk) begin: initialize_ppmatrix
//     if(rst) begin
//         for(int i = 0; i < 64; i++) begin
//             pp[i] <= '0;
//         end
//     end
//     else if(i_rdy) begin
//         for(int i = 0; i < 64; i++) begin
//             for(int j = 0; j < 64; j++) begin
//                 pp[i][j] <= A_reg[j] & B_reg[i];
//             end
//         end 
//     end
// end

// always_comb begin: initialize_ppmatrix
//     if(rst) begin
//         for(int i = 0; i < 32; i++) begin
//             pp[i] = '0;
//         end
//     end
//     else begin
//         for(int i = 0; i < 32; i++) begin
//             for(int j = 0; j < 64; j++) begin
//                 pp[i][j] = A_reg[j] & B_reg[i];
//             end
//         end 
//     end
// end

//stage 0 reduction
HA ha0( .a(A_reg[0] & B_reg[28]), .b(A_reg[1] & B_reg[27]), .sum(s0[0]), .cout(c0[0]) );
FA fa0( .a(A_reg[0] & B_reg[29]), .b(A_reg[1] & B_reg[28]), .cin(A_reg[2] & B_reg[27]), .sum(s0[1]), .cout(c0[1]) );
HA ha1( .a(A_reg[4] & B_reg[25]), .b(A_reg[5] & B_reg[24]), .sum(s0[2]), .cout(c0[2]) );
FA fa1( .a(A_reg[0] & B_reg[30]), .b(A_reg[1] & B_reg[29]), .cin(A_reg[2] & B_reg[28]), .sum(s0[3]), .cout(c0[3]) );
FA fa2( .a(A_reg[4] & B_reg[26]), .b(A_reg[5] & B_reg[25]), .cin(A_reg[6] & B_reg[24]), .sum(s0[4]), .cout(c0[4]) );
HA ha2( .a(A_reg[8] & B_reg[22]), .b(A_reg[9] & B_reg[21]), .sum(s0[5]), .cout(c0[5]) );
FA fa3( .a(A_reg[0] & B_reg[31]), .b(A_reg[1] & B_reg[30]), .cin(A_reg[2] & B_reg[29]), .sum(s0[6]), .cout(c0[6]) );
FA fa4( .a(A_reg[4] & B_reg[27]), .b(A_reg[5] & B_reg[26]), .cin(A_reg[6] & B_reg[25]), .sum(s0[7]), .cout(c0[7]) );
FA fa5( .a(A_reg[8] & B_reg[23]), .b(A_reg[9] & B_reg[22]), .cin(A_reg[10] & B_reg[21]), .sum(s0[8]), .cout(c0[8]) );
HA ha3( .a(A_reg[12] & B_reg[19]), .b(A_reg[13] & B_reg[18]), .sum(s0[9]), .cout(c0[9]) );
FA fa6( .a(A_reg[1] & B_reg[31]), .b(A_reg[2] & B_reg[30]), .cin(A_reg[3] & B_reg[29]), .sum(s0[10]), .cout(c0[10]) );
FA fa7( .a(A_reg[5] & B_reg[27]), .b(A_reg[6] & B_reg[26]), .cin(A_reg[7] & B_reg[25]), .sum(s0[11]), .cout(c0[11]) );
FA fa8( .a(A_reg[9] & B_reg[23]), .b(A_reg[10] & B_reg[22]), .cin(A_reg[11] & B_reg[21]), .sum(s0[12]), .cout(c0[12]) );
HA ha4( .a(A_reg[13] & B_reg[19]), .b(A_reg[14] & B_reg[18]), .sum(s0[13]), .cout(c0[13]) );
FA fa9( .a(A_reg[2] & B_reg[31]), .b(A_reg[3] & B_reg[30]), .cin(A_reg[4] & B_reg[29]), .sum(s0[14]), .cout(c0[14]) );
FA fa10( .a(A_reg[6] & B_reg[27]), .b(A_reg[7] & B_reg[26]), .cin(A_reg[8] & B_reg[25]), .sum(s0[15]), .cout(c0[15]) );
FA fa11( .a(A_reg[10] & B_reg[23]), .b(A_reg[11] & B_reg[22]), .cin(A_reg[12] & B_reg[21]), .sum(s0[16]), .cout(c0[16]) );
FA fa12( .a(A_reg[3] & B_reg[31]), .b(A_reg[4] & B_reg[30]), .cin(A_reg[5] & B_reg[29]), .sum(s0[17]), .cout(c0[17]) );
FA fa13( .a(A_reg[7] & B_reg[27]), .b(A_reg[8] & B_reg[26]), .cin(A_reg[9] & B_reg[25]), .sum(s0[18]), .cout(c0[18]) );
FA fa14( .a(A_reg[4] & B_reg[31]), .b(A_reg[5] & B_reg[30]), .cin(A_reg[6] & B_reg[29]), .sum(s0[19]), .cout(c0[19]) );
//stage 1 reduction
HA ha5( .a(A_reg[0] & B_reg[19]), .b(A_reg[1] & B_reg[18]), .sum(s1[0]), .cout(c1[0]) );
FA fa15( .a(A_reg[0] & B_reg[20]), .b(A_reg[1] & B_reg[19]), .cin(A_reg[2] & B_reg[18]), .sum(s1[1]), .cout(c1[1]) );
HA ha6( .a(A_reg[4] & B_reg[16]), .b(A_reg[5] & B_reg[15]), .sum(s1[2]), .cout(c1[2]) );
FA fa16( .a(A_reg[0] & B_reg[21]), .b(A_reg[1] & B_reg[20]), .cin(A_reg[2] & B_reg[19]), .sum(s1[3]), .cout(c1[3]) );
FA fa17( .a(A_reg[4] & B_reg[17]), .b(A_reg[5] & B_reg[16]), .cin(A_reg[6] & B_reg[15]), .sum(s1[4]), .cout(c1[4]) );
HA ha7( .a(A_reg[8] & B_reg[13]), .b(A_reg[9] & B_reg[12]), .sum(s1[5]), .cout(c1[5]) );
FA fa18( .a(A_reg[0] & B_reg[22]), .b(A_reg[1] & B_reg[21]), .cin(A_reg[2] & B_reg[20]), .sum(s1[6]), .cout(c1[6]) );
FA fa19( .a(A_reg[4] & B_reg[18]), .b(A_reg[5] & B_reg[17]), .cin(A_reg[6] & B_reg[16]), .sum(s1[7]), .cout(c1[7]) );
FA fa20( .a(A_reg[8] & B_reg[14]), .b(A_reg[9] & B_reg[13]), .cin(A_reg[10] & B_reg[12]), .sum(s1[8]), .cout(c1[8]) );
HA ha8( .a(A_reg[12] & B_reg[10]), .b(A_reg[13] & B_reg[9]), .sum(s1[9]), .cout(c1[9]) );
FA fa21( .a(A_reg[0] & B_reg[23]), .b(A_reg[1] & B_reg[22]), .cin(A_reg[2] & B_reg[21]), .sum(s1[10]), .cout(c1[10]) );
FA fa22( .a(A_reg[4] & B_reg[19]), .b(A_reg[5] & B_reg[18]), .cin(A_reg[6] & B_reg[17]), .sum(s1[11]), .cout(c1[11]) );
FA fa23( .a(A_reg[8] & B_reg[15]), .b(A_reg[9] & B_reg[14]), .cin(A_reg[10] & B_reg[13]), .sum(s1[12]), .cout(c1[12]) );
FA fa24( .a(A_reg[12] & B_reg[11]), .b(A_reg[13] & B_reg[10]), .cin(A_reg[14] & B_reg[9]), .sum(s1[13]), .cout(c1[13]) );
HA ha9( .a(A_reg[16] & B_reg[7]), .b(A_reg[17] & B_reg[6]), .sum(s1[14]), .cout(c1[14]) );
FA fa25( .a(A_reg[0] & B_reg[24]), .b(A_reg[1] & B_reg[23]), .cin(A_reg[2] & B_reg[22]), .sum(s1[15]), .cout(c1[15]) );
FA fa26( .a(A_reg[4] & B_reg[20]), .b(A_reg[5] & B_reg[19]), .cin(A_reg[6] & B_reg[18]), .sum(s1[16]), .cout(c1[16]) );
FA fa27( .a(A_reg[8] & B_reg[16]), .b(A_reg[9] & B_reg[15]), .cin(A_reg[10] & B_reg[14]), .sum(s1[17]), .cout(c1[17]) );
FA fa28( .a(A_reg[12] & B_reg[12]), .b(A_reg[13] & B_reg[11]), .cin(A_reg[14] & B_reg[10]), .sum(s1[18]), .cout(c1[18]) );
FA fa29( .a(A_reg[16] & B_reg[8]), .b(A_reg[17] & B_reg[7]), .cin(A_reg[18] & B_reg[6]), .sum(s1[19]), .cout(c1[19]) );
HA ha10( .a(A_reg[20] & B_reg[4]), .b(A_reg[21] & B_reg[3]), .sum(s1[20]), .cout(c1[20]) );
FA fa30( .a(A_reg[0] & B_reg[25]), .b(A_reg[1] & B_reg[24]), .cin(A_reg[2] & B_reg[23]), .sum(s1[21]), .cout(c1[21]) );
FA fa31( .a(A_reg[4] & B_reg[21]), .b(A_reg[5] & B_reg[20]), .cin(A_reg[6] & B_reg[19]), .sum(s1[22]), .cout(c1[22]) );
FA fa32( .a(A_reg[8] & B_reg[17]), .b(A_reg[9] & B_reg[16]), .cin(A_reg[10] & B_reg[15]), .sum(s1[23]), .cout(c1[23]) );
FA fa33( .a(A_reg[12] & B_reg[13]), .b(A_reg[13] & B_reg[12]), .cin(A_reg[14] & B_reg[11]), .sum(s1[24]), .cout(c1[24]) );
FA fa34( .a(A_reg[16] & B_reg[9]), .b(A_reg[17] & B_reg[8]), .cin(A_reg[18] & B_reg[7]), .sum(s1[25]), .cout(c1[25]) );
FA fa35( .a(A_reg[20] & B_reg[5]), .b(A_reg[21] & B_reg[4]), .cin(A_reg[22] & B_reg[3]), .sum(s1[26]), .cout(c1[26]) );
HA ha11( .a(A_reg[24] & B_reg[1]), .b(A_reg[25] & B_reg[0]), .sum(s1[27]), .cout(c1[27]) );
FA fa36( .a(A_reg[0] & B_reg[26]), .b(A_reg[1] & B_reg[25]), .cin(A_reg[2] & B_reg[24]), .sum(s1[28]), .cout(c1[28]) );
FA fa37( .a(A_reg[4] & B_reg[22]), .b(A_reg[5] & B_reg[21]), .cin(A_reg[6] & B_reg[20]), .sum(s1[29]), .cout(c1[29]) );
FA fa38( .a(A_reg[8] & B_reg[18]), .b(A_reg[9] & B_reg[17]), .cin(A_reg[10] & B_reg[16]), .sum(s1[30]), .cout(c1[30]) );
FA fa39( .a(A_reg[12] & B_reg[14]), .b(A_reg[13] & B_reg[13]), .cin(A_reg[14] & B_reg[12]), .sum(s1[31]), .cout(c1[31]) );
FA fa40( .a(A_reg[16] & B_reg[10]), .b(A_reg[17] & B_reg[9]), .cin(A_reg[18] & B_reg[8]), .sum(s1[32]), .cout(c1[32]) );
FA fa41( .a(A_reg[20] & B_reg[6]), .b(A_reg[21] & B_reg[5]), .cin(A_reg[22] & B_reg[4]), .sum(s1[33]), .cout(c1[33]) );
FA fa42( .a(A_reg[24] & B_reg[2]), .b(A_reg[25] & B_reg[1]), .cin(A_reg[26] & B_reg[0]), .sum(s1[34]), .cout(c1[34]) );
HA ha12( .a(c1[22]), .b(c1[23]), .sum(s1[35]), .cout(c1[35]) );
FA fa43( .a(A_reg[0] & B_reg[27]), .b(A_reg[1] & B_reg[26]), .cin(A_reg[2] & B_reg[25]), .sum(s1[36]), .cout(c1[36]) );
FA fa44( .a(A_reg[4] & B_reg[23]), .b(A_reg[5] & B_reg[22]), .cin(A_reg[6] & B_reg[21]), .sum(s1[37]), .cout(c1[37]) );
FA fa45( .a(A_reg[8] & B_reg[19]), .b(A_reg[9] & B_reg[18]), .cin(A_reg[10] & B_reg[17]), .sum(s1[38]), .cout(c1[38]) );
FA fa46( .a(A_reg[12] & B_reg[15]), .b(A_reg[13] & B_reg[14]), .cin(A_reg[14] & B_reg[13]), .sum(s1[39]), .cout(c1[39]) );
FA fa47( .a(A_reg[16] & B_reg[11]), .b(A_reg[17] & B_reg[10]), .cin(A_reg[18] & B_reg[9]), .sum(s1[40]), .cout(c1[40]) );
FA fa48( .a(A_reg[20] & B_reg[7]), .b(A_reg[21] & B_reg[6]), .cin(A_reg[22] & B_reg[5]), .sum(s1[41]), .cout(c1[41]) );
FA fa49( .a(A_reg[24] & B_reg[3]), .b(A_reg[25] & B_reg[2]), .cin(A_reg[26] & B_reg[1]), .sum(s1[42]), .cout(c1[42]) );
FA fa50( .a(c1[28]), .b(c1[29]), .cin(c1[30]), .sum(s1[43]), .cout(c1[43]) );
HA ha13( .a(c1[32]), .b(c1[33]), .sum(s1[44]), .cout(c1[44]) );
FA fa51( .a(A_reg[2] & B_reg[26]), .b(A_reg[3] & B_reg[25]), .cin(A_reg[4] & B_reg[24]), .sum(s1[45]), .cout(c1[45]) );
FA fa52( .a(A_reg[6] & B_reg[22]), .b(A_reg[7] & B_reg[21]), .cin(A_reg[8] & B_reg[20]), .sum(s1[46]), .cout(c1[46]) );
FA fa53( .a(A_reg[10] & B_reg[18]), .b(A_reg[11] & B_reg[17]), .cin(A_reg[12] & B_reg[16]), .sum(s1[47]), .cout(c1[47]) );
FA fa54( .a(A_reg[14] & B_reg[14]), .b(A_reg[15] & B_reg[13]), .cin(A_reg[16] & B_reg[12]), .sum(s1[48]), .cout(c1[48]) );
FA fa55( .a(A_reg[18] & B_reg[10]), .b(A_reg[19] & B_reg[9]), .cin(A_reg[20] & B_reg[8]), .sum(s1[49]), .cout(c1[49]) );
FA fa56( .a(A_reg[22] & B_reg[6]), .b(A_reg[23] & B_reg[5]), .cin(A_reg[24] & B_reg[4]), .sum(s1[50]), .cout(c1[50]) );
FA fa57( .a(A_reg[26] & B_reg[2]), .b(A_reg[27] & B_reg[1]), .cin(A_reg[28] & B_reg[0]), .sum(s1[51]), .cout(c1[51]) );
FA fa58( .a(c1[36]), .b(c1[37]), .cin(c1[38]), .sum(s1[52]), .cout(c1[52]) );
FA fa59( .a(c1[40]), .b(c1[41]), .cin(c1[42]), .sum(s1[53]), .cout(c1[53]) );
FA fa60( .a(A_reg[3] & B_reg[26]), .b(A_reg[6] & B_reg[23]), .cin(A_reg[7] & B_reg[22]), .sum(s1[54]), .cout(c1[54]) );
FA fa61( .a(A_reg[9] & B_reg[20]), .b(A_reg[10] & B_reg[19]), .cin(A_reg[11] & B_reg[18]), .sum(s1[55]), .cout(c1[55]) );
FA fa62( .a(A_reg[13] & B_reg[16]), .b(A_reg[14] & B_reg[15]), .cin(A_reg[15] & B_reg[14]), .sum(s1[56]), .cout(c1[56]) );
FA fa63( .a(A_reg[17] & B_reg[12]), .b(A_reg[18] & B_reg[11]), .cin(A_reg[19] & B_reg[10]), .sum(s1[57]), .cout(c1[57]) );
FA fa64( .a(A_reg[21] & B_reg[8]), .b(A_reg[22] & B_reg[7]), .cin(A_reg[23] & B_reg[6]), .sum(s1[58]), .cout(c1[58]) );
FA fa65( .a(A_reg[25] & B_reg[4]), .b(A_reg[26] & B_reg[3]), .cin(A_reg[27] & B_reg[2]), .sum(s1[59]), .cout(c1[59]) );
FA fa66( .a(A_reg[29] & B_reg[0]), .b(c0[0]), .cin(s0[1]), .sum(s1[60]), .cout(c1[60]) );
FA fa67( .a(c1[45]), .b(c1[46]), .cin(c1[47]), .sum(s1[61]), .cout(c1[61]) );
FA fa68( .a(c1[49]), .b(c1[50]), .cin(c1[51]), .sum(s1[62]), .cout(c1[62]) );
FA fa69( .a(A_reg[3] & B_reg[27]), .b(A_reg[7] & B_reg[23]), .cin(A_reg[10] & B_reg[20]), .sum(s1[63]), .cout(c1[63]) );
FA fa70( .a(A_reg[12] & B_reg[18]), .b(A_reg[13] & B_reg[17]), .cin(A_reg[14] & B_reg[16]), .sum(s1[64]), .cout(c1[64]) );
FA fa71( .a(A_reg[16] & B_reg[14]), .b(A_reg[17] & B_reg[13]), .cin(A_reg[18] & B_reg[12]), .sum(s1[65]), .cout(c1[65]) );
FA fa72( .a(A_reg[20] & B_reg[10]), .b(A_reg[21] & B_reg[9]), .cin(A_reg[22] & B_reg[8]), .sum(s1[66]), .cout(c1[66]) );
FA fa73( .a(A_reg[24] & B_reg[6]), .b(A_reg[25] & B_reg[5]), .cin(A_reg[26] & B_reg[4]), .sum(s1[67]), .cout(c1[67]) );
FA fa74( .a(A_reg[28] & B_reg[2]), .b(A_reg[29] & B_reg[1]), .cin(A_reg[30] & B_reg[0]), .sum(s1[68]), .cout(c1[68]) );
FA fa75( .a(c0[2]), .b(s0[3]), .cin(s0[4]), .sum(s1[69]), .cout(c1[69]) );
FA fa76( .a(c1[54]), .b(c1[55]), .cin(c1[56]), .sum(s1[70]), .cout(c1[70]) );
FA fa77( .a(c1[58]), .b(c1[59]), .cin(c1[60]), .sum(s1[71]), .cout(c1[71]) );
FA fa78( .a(A_reg[3] & B_reg[28]), .b(A_reg[7] & B_reg[24]), .cin(A_reg[11] & B_reg[20]), .sum(s1[72]), .cout(c1[72]) );
FA fa79( .a(A_reg[15] & B_reg[16]), .b(A_reg[16] & B_reg[15]), .cin(A_reg[17] & B_reg[14]), .sum(s1[73]), .cout(c1[73]) );
FA fa80( .a(A_reg[19] & B_reg[12]), .b(A_reg[20] & B_reg[11]), .cin(A_reg[21] & B_reg[10]), .sum(s1[74]), .cout(c1[74]) );
FA fa81( .a(A_reg[23] & B_reg[8]), .b(A_reg[24] & B_reg[7]), .cin(A_reg[25] & B_reg[6]), .sum(s1[75]), .cout(c1[75]) );
FA fa82( .a(A_reg[27] & B_reg[4]), .b(A_reg[28] & B_reg[3]), .cin(A_reg[29] & B_reg[2]), .sum(s1[76]), .cout(c1[76]) );
FA fa83( .a(A_reg[31] & B_reg[0]), .b(c0[3]), .cin(c0[4]), .sum(s1[77]), .cout(c1[77]) );
FA fa84( .a(s0[6]), .b(s0[7]), .cin(s0[8]), .sum(s1[78]), .cout(c1[78]) );
FA fa85( .a(c1[63]), .b(c1[64]), .cin(c1[65]), .sum(s1[79]), .cout(c1[79]) );
FA fa86( .a(c1[67]), .b(c1[68]), .cin(c1[69]), .sum(s1[80]), .cout(c1[80]) );
FA fa87( .a(A_reg[4] & B_reg[28]), .b(A_reg[8] & B_reg[24]), .cin(A_reg[12] & B_reg[20]), .sum(s1[81]), .cout(c1[81]) );
FA fa88( .a(A_reg[16] & B_reg[16]), .b(A_reg[17] & B_reg[15]), .cin(A_reg[18] & B_reg[14]), .sum(s1[82]), .cout(c1[82]) );
FA fa89( .a(A_reg[20] & B_reg[12]), .b(A_reg[21] & B_reg[11]), .cin(A_reg[22] & B_reg[10]), .sum(s1[83]), .cout(c1[83]) );
FA fa90( .a(A_reg[24] & B_reg[8]), .b(A_reg[25] & B_reg[7]), .cin(A_reg[26] & B_reg[6]), .sum(s1[84]), .cout(c1[84]) );
FA fa91( .a(A_reg[28] & B_reg[4]), .b(A_reg[29] & B_reg[3]), .cin(A_reg[30] & B_reg[2]), .sum(s1[85]), .cout(c1[85]) );
FA fa92( .a(c0[6]), .b(c0[7]), .cin(c0[8]), .sum(s1[86]), .cout(c1[86]) );
FA fa93( .a(s0[10]), .b(s0[11]), .cin(s0[12]), .sum(s1[87]), .cout(c1[87]) );
FA fa94( .a(c1[72]), .b(c1[73]), .cin(c1[74]), .sum(s1[88]), .cout(c1[88]) );
FA fa95( .a(c1[76]), .b(c1[77]), .cin(c1[78]), .sum(s1[89]), .cout(c1[89]) );
FA fa96( .a(A_reg[5] & B_reg[28]), .b(A_reg[9] & B_reg[24]), .cin(A_reg[13] & B_reg[20]), .sum(s1[90]), .cout(c1[90]) );
FA fa97( .a(A_reg[15] & B_reg[18]), .b(A_reg[16] & B_reg[17]), .cin(A_reg[17] & B_reg[16]), .sum(s1[91]), .cout(c1[91]) );
FA fa98( .a(A_reg[19] & B_reg[14]), .b(A_reg[20] & B_reg[13]), .cin(A_reg[21] & B_reg[12]), .sum(s1[92]), .cout(c1[92]) );
FA fa99( .a(A_reg[23] & B_reg[10]), .b(A_reg[24] & B_reg[9]), .cin(A_reg[25] & B_reg[8]), .sum(s1[93]), .cout(c1[93]) );
FA fa100( .a(A_reg[27] & B_reg[6]), .b(A_reg[28] & B_reg[5]), .cin(A_reg[29] & B_reg[4]), .sum(s1[94]), .cout(c1[94]) );
FA fa101( .a(A_reg[31] & B_reg[2]), .b(c0[10]), .cin(c0[11]), .sum(s1[95]), .cout(c1[95]) );
FA fa102( .a(c0[13]), .b(s0[14]), .cin(s0[15]), .sum(s1[96]), .cout(c1[96]) );
FA fa103( .a(c1[81]), .b(c1[82]), .cin(c1[83]), .sum(s1[97]), .cout(c1[97]) );
FA fa104( .a(c1[85]), .b(c1[86]), .cin(c1[87]), .sum(s1[98]), .cout(c1[98]) );
FA fa105( .a(A_reg[6] & B_reg[28]), .b(A_reg[10] & B_reg[24]), .cin(A_reg[11] & B_reg[23]), .sum(s1[99]), .cout(c1[99]) );
FA fa106( .a(A_reg[13] & B_reg[21]), .b(A_reg[14] & B_reg[20]), .cin(A_reg[15] & B_reg[19]), .sum(s1[100]), .cout(c1[100]) );
FA fa107( .a(A_reg[17] & B_reg[17]), .b(A_reg[18] & B_reg[16]), .cin(A_reg[19] & B_reg[15]), .sum(s1[101]), .cout(c1[101]) );
FA fa108( .a(A_reg[21] & B_reg[13]), .b(A_reg[22] & B_reg[12]), .cin(A_reg[23] & B_reg[11]), .sum(s1[102]), .cout(c1[102]) );
FA fa109( .a(A_reg[25] & B_reg[9]), .b(A_reg[26] & B_reg[8]), .cin(A_reg[27] & B_reg[7]), .sum(s1[103]), .cout(c1[103]) );
FA fa110( .a(A_reg[29] & B_reg[5]), .b(A_reg[30] & B_reg[4]), .cin(A_reg[31] & B_reg[3]), .sum(s1[104]), .cout(c1[104]) );
FA fa111( .a(c0[15]), .b(c0[16]), .cin(s0[17]), .sum(s1[105]), .cout(c1[105]) );
FA fa112( .a(c1[90]), .b(c1[91]), .cin(c1[92]), .sum(s1[106]), .cout(c1[106]) );
FA fa113( .a(c1[94]), .b(c1[95]), .cin(c1[96]), .sum(s1[107]), .cout(c1[107]) );
FA fa114( .a(A_reg[7] & B_reg[28]), .b(A_reg[8] & B_reg[27]), .cin(A_reg[9] & B_reg[26]), .sum(s1[108]), .cout(c1[108]) );
FA fa115( .a(A_reg[11] & B_reg[24]), .b(A_reg[12] & B_reg[23]), .cin(A_reg[13] & B_reg[22]), .sum(s1[109]), .cout(c1[109]) );
FA fa116( .a(A_reg[15] & B_reg[20]), .b(A_reg[16] & B_reg[19]), .cin(A_reg[17] & B_reg[18]), .sum(s1[110]), .cout(c1[110]) );
FA fa117( .a(A_reg[19] & B_reg[16]), .b(A_reg[20] & B_reg[15]), .cin(A_reg[21] & B_reg[14]), .sum(s1[111]), .cout(c1[111]) );
FA fa118( .a(A_reg[23] & B_reg[12]), .b(A_reg[24] & B_reg[11]), .cin(A_reg[25] & B_reg[10]), .sum(s1[112]), .cout(c1[112]) );
FA fa119( .a(A_reg[27] & B_reg[8]), .b(A_reg[28] & B_reg[7]), .cin(A_reg[29] & B_reg[6]), .sum(s1[113]), .cout(c1[113]) );
FA fa120( .a(A_reg[31] & B_reg[4]), .b(c0[17]), .cin(c0[18]), .sum(s1[114]), .cout(c1[114]) );
FA fa121( .a(c1[99]), .b(c1[100]), .cin(c1[101]), .sum(s1[115]), .cout(c1[115]) );
FA fa122( .a(c1[103]), .b(c1[104]), .cin(c1[105]), .sum(s1[116]), .cout(c1[116]) );
FA fa123( .a(A_reg[5] & B_reg[31]), .b(A_reg[6] & B_reg[30]), .cin(A_reg[7] & B_reg[29]), .sum(s1[117]), .cout(c1[117]) );
FA fa124( .a(A_reg[9] & B_reg[27]), .b(A_reg[10] & B_reg[26]), .cin(A_reg[11] & B_reg[25]), .sum(s1[118]), .cout(c1[118]) );
FA fa125( .a(A_reg[13] & B_reg[23]), .b(A_reg[14] & B_reg[22]), .cin(A_reg[15] & B_reg[21]), .sum(s1[119]), .cout(c1[119]) );
FA fa126( .a(A_reg[17] & B_reg[19]), .b(A_reg[18] & B_reg[18]), .cin(A_reg[19] & B_reg[17]), .sum(s1[120]), .cout(c1[120]) );
FA fa127( .a(A_reg[21] & B_reg[15]), .b(A_reg[22] & B_reg[14]), .cin(A_reg[23] & B_reg[13]), .sum(s1[121]), .cout(c1[121]) );
FA fa128( .a(A_reg[25] & B_reg[11]), .b(A_reg[26] & B_reg[10]), .cin(A_reg[27] & B_reg[9]), .sum(s1[122]), .cout(c1[122]) );
FA fa129( .a(A_reg[29] & B_reg[7]), .b(A_reg[30] & B_reg[6]), .cin(A_reg[31] & B_reg[5]), .sum(s1[123]), .cout(c1[123]) );
FA fa130( .a(c1[108]), .b(c1[109]), .cin(c1[110]), .sum(s1[124]), .cout(c1[124]) );
FA fa131( .a(c1[112]), .b(c1[113]), .cin(c1[114]), .sum(s1[125]), .cout(c1[125]) );
FA fa132( .a(A_reg[6] & B_reg[31]), .b(A_reg[7] & B_reg[30]), .cin(A_reg[8] & B_reg[29]), .sum(s1[126]), .cout(c1[126]) );
FA fa133( .a(A_reg[10] & B_reg[27]), .b(A_reg[11] & B_reg[26]), .cin(A_reg[12] & B_reg[25]), .sum(s1[127]), .cout(c1[127]) );
FA fa134( .a(A_reg[14] & B_reg[23]), .b(A_reg[15] & B_reg[22]), .cin(A_reg[16] & B_reg[21]), .sum(s1[128]), .cout(c1[128]) );
FA fa135( .a(A_reg[18] & B_reg[19]), .b(A_reg[19] & B_reg[18]), .cin(A_reg[20] & B_reg[17]), .sum(s1[129]), .cout(c1[129]) );
FA fa136( .a(A_reg[22] & B_reg[15]), .b(A_reg[23] & B_reg[14]), .cin(A_reg[24] & B_reg[13]), .sum(s1[130]), .cout(c1[130]) );
FA fa137( .a(A_reg[26] & B_reg[11]), .b(A_reg[27] & B_reg[10]), .cin(A_reg[28] & B_reg[9]), .sum(s1[131]), .cout(c1[131]) );
FA fa138( .a(A_reg[30] & B_reg[7]), .b(A_reg[31] & B_reg[6]), .cin(c1[117]), .sum(s1[132]), .cout(c1[132]) );
FA fa139( .a(c1[119]), .b(c1[120]), .cin(c1[121]), .sum(s1[133]), .cout(c1[133]) );
FA fa140( .a(A_reg[7] & B_reg[31]), .b(A_reg[8] & B_reg[30]), .cin(A_reg[9] & B_reg[29]), .sum(s1[134]), .cout(c1[134]) );
FA fa141( .a(A_reg[11] & B_reg[27]), .b(A_reg[12] & B_reg[26]), .cin(A_reg[13] & B_reg[25]), .sum(s1[135]), .cout(c1[135]) );
FA fa142( .a(A_reg[15] & B_reg[23]), .b(A_reg[16] & B_reg[22]), .cin(A_reg[17] & B_reg[21]), .sum(s1[136]), .cout(c1[136]) );
FA fa143( .a(A_reg[19] & B_reg[19]), .b(A_reg[20] & B_reg[18]), .cin(A_reg[21] & B_reg[17]), .sum(s1[137]), .cout(c1[137]) );
FA fa144( .a(A_reg[23] & B_reg[15]), .b(A_reg[24] & B_reg[14]), .cin(A_reg[25] & B_reg[13]), .sum(s1[138]), .cout(c1[138]) );
FA fa145( .a(A_reg[27] & B_reg[11]), .b(A_reg[28] & B_reg[10]), .cin(A_reg[29] & B_reg[9]), .sum(s1[139]), .cout(c1[139]) );
FA fa146( .a(A_reg[31] & B_reg[7]), .b(c1[126]), .cin(c1[127]), .sum(s1[140]), .cout(c1[140]) );
FA fa147( .a(A_reg[8] & B_reg[31]), .b(A_reg[9] & B_reg[30]), .cin(A_reg[10] & B_reg[29]), .sum(s1[141]), .cout(c1[141]) );
FA fa148( .a(A_reg[12] & B_reg[27]), .b(A_reg[13] & B_reg[26]), .cin(A_reg[14] & B_reg[25]), .sum(s1[142]), .cout(c1[142]) );
FA fa149( .a(A_reg[16] & B_reg[23]), .b(A_reg[17] & B_reg[22]), .cin(A_reg[18] & B_reg[21]), .sum(s1[143]), .cout(c1[143]) );
FA fa150( .a(A_reg[20] & B_reg[19]), .b(A_reg[21] & B_reg[18]), .cin(A_reg[22] & B_reg[17]), .sum(s1[144]), .cout(c1[144]) );
FA fa151( .a(A_reg[24] & B_reg[15]), .b(A_reg[25] & B_reg[14]), .cin(A_reg[26] & B_reg[13]), .sum(s1[145]), .cout(c1[145]) );
FA fa152( .a(A_reg[28] & B_reg[11]), .b(A_reg[29] & B_reg[10]), .cin(A_reg[30] & B_reg[9]), .sum(s1[146]), .cout(c1[146]) );
FA fa153( .a(A_reg[9] & B_reg[31]), .b(A_reg[10] & B_reg[30]), .cin(A_reg[11] & B_reg[29]), .sum(s1[147]), .cout(c1[147]) );
FA fa154( .a(A_reg[13] & B_reg[27]), .b(A_reg[14] & B_reg[26]), .cin(A_reg[15] & B_reg[25]), .sum(s1[148]), .cout(c1[148]) );
FA fa155( .a(A_reg[17] & B_reg[23]), .b(A_reg[18] & B_reg[22]), .cin(A_reg[19] & B_reg[21]), .sum(s1[149]), .cout(c1[149]) );
FA fa156( .a(A_reg[21] & B_reg[19]), .b(A_reg[22] & B_reg[18]), .cin(A_reg[23] & B_reg[17]), .sum(s1[150]), .cout(c1[150]) );
FA fa157( .a(A_reg[25] & B_reg[15]), .b(A_reg[26] & B_reg[14]), .cin(A_reg[27] & B_reg[13]), .sum(s1[151]), .cout(c1[151]) );
FA fa158( .a(A_reg[10] & B_reg[31]), .b(A_reg[11] & B_reg[30]), .cin(A_reg[12] & B_reg[29]), .sum(s1[152]), .cout(c1[152]) );
FA fa159( .a(A_reg[14] & B_reg[27]), .b(A_reg[15] & B_reg[26]), .cin(A_reg[16] & B_reg[25]), .sum(s1[153]), .cout(c1[153]) );
FA fa160( .a(A_reg[18] & B_reg[23]), .b(A_reg[19] & B_reg[22]), .cin(A_reg[20] & B_reg[21]), .sum(s1[154]), .cout(c1[154]) );
FA fa161( .a(A_reg[22] & B_reg[19]), .b(A_reg[23] & B_reg[18]), .cin(A_reg[24] & B_reg[17]), .sum(s1[155]), .cout(c1[155]) );
FA fa162( .a(A_reg[11] & B_reg[31]), .b(A_reg[12] & B_reg[30]), .cin(A_reg[13] & B_reg[29]), .sum(s1[156]), .cout(c1[156]) );
FA fa163( .a(A_reg[15] & B_reg[27]), .b(A_reg[16] & B_reg[26]), .cin(A_reg[17] & B_reg[25]), .sum(s1[157]), .cout(c1[157]) );
FA fa164( .a(A_reg[19] & B_reg[23]), .b(A_reg[20] & B_reg[22]), .cin(A_reg[21] & B_reg[21]), .sum(s1[158]), .cout(c1[158]) );
FA fa165( .a(A_reg[12] & B_reg[31]), .b(A_reg[13] & B_reg[30]), .cin(A_reg[14] & B_reg[29]), .sum(s1[159]), .cout(c1[159]) );
FA fa166( .a(A_reg[16] & B_reg[27]), .b(A_reg[17] & B_reg[26]), .cin(A_reg[18] & B_reg[25]), .sum(s1[160]), .cout(c1[160]) );
FA fa167( .a(A_reg[13] & B_reg[31]), .b(A_reg[14] & B_reg[30]), .cin(A_reg[15] & B_reg[29]), .sum(s1[161]), .cout(c1[161]) );
//stage 2 reduction
HA ha14( .a(A_reg[0] & B_reg[13]), .b(A_reg[1] & B_reg[12]), .sum(s2[0]), .cout(c2[0]) );
FA fa168( .a(A_reg[0] & B_reg[14]), .b(A_reg[1] & B_reg[13]), .cin(A_reg[2] & B_reg[12]), .sum(s2[1]), .cout(c2[1]) );
HA ha15( .a(A_reg[4] & B_reg[10]), .b(A_reg[5] & B_reg[9]), .sum(s2[2]), .cout(c2[2]) );
FA fa169( .a(A_reg[0] & B_reg[15]), .b(A_reg[1] & B_reg[14]), .cin(A_reg[2] & B_reg[13]), .sum(s2[3]), .cout(c2[3]) );
FA fa170( .a(A_reg[4] & B_reg[11]), .b(A_reg[5] & B_reg[10]), .cin(A_reg[6] & B_reg[9]), .sum(s2[4]), .cout(c2[4]) );
HA ha16( .a(A_reg[8] & B_reg[7]), .b(A_reg[9] & B_reg[6]), .sum(s2[5]), .cout(c2[5]) );
FA fa171( .a(A_reg[0] & B_reg[16]), .b(A_reg[1] & B_reg[15]), .cin(A_reg[2] & B_reg[14]), .sum(s2[6]), .cout(c2[6]) );
FA fa172( .a(A_reg[4] & B_reg[12]), .b(A_reg[5] & B_reg[11]), .cin(A_reg[6] & B_reg[10]), .sum(s2[7]), .cout(c2[7]) );
FA fa173( .a(A_reg[8] & B_reg[8]), .b(A_reg[9] & B_reg[7]), .cin(A_reg[10] & B_reg[6]), .sum(s2[8]), .cout(c2[8]) );
HA ha17( .a(A_reg[12] & B_reg[4]), .b(A_reg[13] & B_reg[3]), .sum(s2[9]), .cout(c2[9]) );
FA fa174( .a(A_reg[0] & B_reg[17]), .b(A_reg[1] & B_reg[16]), .cin(A_reg[2] & B_reg[15]), .sum(s2[10]), .cout(c2[10]) );
FA fa175( .a(A_reg[4] & B_reg[13]), .b(A_reg[5] & B_reg[12]), .cin(A_reg[6] & B_reg[11]), .sum(s2[11]), .cout(c2[11]) );
FA fa176( .a(A_reg[8] & B_reg[9]), .b(A_reg[9] & B_reg[8]), .cin(A_reg[10] & B_reg[7]), .sum(s2[12]), .cout(c2[12]) );
FA fa177( .a(A_reg[12] & B_reg[5]), .b(A_reg[13] & B_reg[4]), .cin(A_reg[14] & B_reg[3]), .sum(s2[13]), .cout(c2[13]) );
HA ha18( .a(A_reg[16] & B_reg[1]), .b(A_reg[17] & B_reg[0]), .sum(s2[14]), .cout(c2[14]) );
FA fa178( .a(A_reg[0] & B_reg[18]), .b(A_reg[1] & B_reg[17]), .cin(A_reg[2] & B_reg[16]), .sum(s2[15]), .cout(c2[15]) );
FA fa179( .a(A_reg[4] & B_reg[14]), .b(A_reg[5] & B_reg[13]), .cin(A_reg[6] & B_reg[12]), .sum(s2[16]), .cout(c2[16]) );
FA fa180( .a(A_reg[8] & B_reg[10]), .b(A_reg[9] & B_reg[9]), .cin(A_reg[10] & B_reg[8]), .sum(s2[17]), .cout(c2[17]) );
FA fa181( .a(A_reg[12] & B_reg[6]), .b(A_reg[13] & B_reg[5]), .cin(A_reg[14] & B_reg[4]), .sum(s2[18]), .cout(c2[18]) );
FA fa182( .a(A_reg[16] & B_reg[2]), .b(A_reg[17] & B_reg[1]), .cin(A_reg[18] & B_reg[0]), .sum(s2[19]), .cout(c2[19]) );
HA ha19( .a(c2[11]), .b(c2[12]), .sum(s2[20]), .cout(c2[20]) );
FA fa183( .a(A_reg[2] & B_reg[17]), .b(A_reg[3] & B_reg[16]), .cin(A_reg[4] & B_reg[15]), .sum(s2[21]), .cout(c2[21]) );
FA fa184( .a(A_reg[6] & B_reg[13]), .b(A_reg[7] & B_reg[12]), .cin(A_reg[8] & B_reg[11]), .sum(s2[22]), .cout(c2[22]) );
FA fa185( .a(A_reg[10] & B_reg[9]), .b(A_reg[11] & B_reg[8]), .cin(A_reg[12] & B_reg[7]), .sum(s2[23]), .cout(c2[23]) );
FA fa186( .a(A_reg[14] & B_reg[5]), .b(A_reg[15] & B_reg[4]), .cin(A_reg[16] & B_reg[3]), .sum(s2[24]), .cout(c2[24]) );
FA fa187( .a(A_reg[18] & B_reg[1]), .b(A_reg[19] & B_reg[0]), .cin(s1[0]), .sum(s2[25]), .cout(c2[25]) );
FA fa188( .a(c2[16]), .b(c2[17]), .cin(c2[18]), .sum(s2[26]), .cout(c2[26]) );
FA fa189( .a(A_reg[3] & B_reg[17]), .b(A_reg[6] & B_reg[14]), .cin(A_reg[7] & B_reg[13]), .sum(s2[27]), .cout(c2[27]) );
FA fa190( .a(A_reg[9] & B_reg[11]), .b(A_reg[10] & B_reg[10]), .cin(A_reg[11] & B_reg[9]), .sum(s2[28]), .cout(c2[28]) );
FA fa191( .a(A_reg[13] & B_reg[7]), .b(A_reg[14] & B_reg[6]), .cin(A_reg[15] & B_reg[5]), .sum(s2[29]), .cout(c2[29]) );
FA fa192( .a(A_reg[17] & B_reg[3]), .b(A_reg[18] & B_reg[2]), .cin(A_reg[19] & B_reg[1]), .sum(s2[30]), .cout(c2[30]) );
FA fa193( .a(c1[0]), .b(s1[1]), .cin(s1[2]), .sum(s2[31]), .cout(c2[31]) );
FA fa194( .a(c2[22]), .b(c2[23]), .cin(c2[24]), .sum(s2[32]), .cout(c2[32]) );
FA fa195( .a(A_reg[3] & B_reg[18]), .b(A_reg[7] & B_reg[14]), .cin(A_reg[10] & B_reg[11]), .sum(s2[33]), .cout(c2[33]) );
FA fa196( .a(A_reg[12] & B_reg[9]), .b(A_reg[13] & B_reg[8]), .cin(A_reg[14] & B_reg[7]), .sum(s2[34]), .cout(c2[34]) );
FA fa197( .a(A_reg[16] & B_reg[5]), .b(A_reg[17] & B_reg[4]), .cin(A_reg[18] & B_reg[3]), .sum(s2[35]), .cout(c2[35]) );
FA fa198( .a(A_reg[20] & B_reg[1]), .b(A_reg[21] & B_reg[0]), .cin(c1[1]), .sum(s2[36]), .cout(c2[36]) );
FA fa199( .a(s1[3]), .b(s1[4]), .cin(s1[5]), .sum(s2[37]), .cout(c2[37]) );
FA fa200( .a(c2[28]), .b(c2[29]), .cin(c2[30]), .sum(s2[38]), .cout(c2[38]) );
FA fa201( .a(A_reg[3] & B_reg[19]), .b(A_reg[7] & B_reg[15]), .cin(A_reg[11] & B_reg[11]), .sum(s2[39]), .cout(c2[39]) );
FA fa202( .a(A_reg[15] & B_reg[7]), .b(A_reg[16] & B_reg[6]), .cin(A_reg[17] & B_reg[5]), .sum(s2[40]), .cout(c2[40]) );
FA fa203( .a(A_reg[19] & B_reg[3]), .b(A_reg[20] & B_reg[2]), .cin(A_reg[21] & B_reg[1]), .sum(s2[41]), .cout(c2[41]) );
FA fa204( .a(c1[3]), .b(c1[4]), .cin(c1[5]), .sum(s2[42]), .cout(c2[42]) );
FA fa205( .a(s1[7]), .b(s1[8]), .cin(s1[9]), .sum(s2[43]), .cout(c2[43]) );
FA fa206( .a(c2[34]), .b(c2[35]), .cin(c2[36]), .sum(s2[44]), .cout(c2[44]) );
FA fa207( .a(A_reg[3] & B_reg[20]), .b(A_reg[7] & B_reg[16]), .cin(A_reg[11] & B_reg[12]), .sum(s2[45]), .cout(c2[45]) );
FA fa208( .a(A_reg[18] & B_reg[5]), .b(A_reg[19] & B_reg[4]), .cin(A_reg[20] & B_reg[3]), .sum(s2[46]), .cout(c2[46]) );
FA fa209( .a(A_reg[22] & B_reg[1]), .b(A_reg[23] & B_reg[0]), .cin(c1[6]), .sum(s2[47]), .cout(c2[47]) );
FA fa210( .a(c1[8]), .b(c1[9]), .cin(s1[10]), .sum(s2[48]), .cout(c2[48]) );
FA fa211( .a(s1[12]), .b(s1[13]), .cin(s1[14]), .sum(s2[49]), .cout(c2[49]) );
FA fa212( .a(c2[40]), .b(c2[41]), .cin(c2[42]), .sum(s2[50]), .cout(c2[50]) );
FA fa213( .a(A_reg[3] & B_reg[21]), .b(A_reg[7] & B_reg[17]), .cin(A_reg[11] & B_reg[13]), .sum(s2[51]), .cout(c2[51]) );
FA fa214( .a(A_reg[19] & B_reg[5]), .b(A_reg[22] & B_reg[2]), .cin(A_reg[23] & B_reg[1]), .sum(s2[52]), .cout(c2[52]) );
FA fa215( .a(c1[10]), .b(c1[11]), .cin(c1[12]), .sum(s2[53]), .cout(c2[53]) );
FA fa216( .a(c1[14]), .b(s1[15]), .cin(s1[16]), .sum(s2[54]), .cout(c2[54]) );
FA fa217( .a(s1[18]), .b(s1[19]), .cin(s1[20]), .sum(s2[55]), .cout(c2[55]) );
FA fa218( .a(c2[46]), .b(c2[47]), .cin(c2[48]), .sum(s2[56]), .cout(c2[56]) );
FA fa219( .a(A_reg[3] & B_reg[22]), .b(A_reg[7] & B_reg[18]), .cin(A_reg[11] & B_reg[14]), .sum(s2[57]), .cout(c2[57]) );
FA fa220( .a(A_reg[19] & B_reg[6]), .b(A_reg[23] & B_reg[2]), .cin(c1[15]), .sum(s2[58]), .cout(c2[58]) );
FA fa221( .a(c1[17]), .b(c1[18]), .cin(c1[19]), .sum(s2[59]), .cout(c2[59]) );
FA fa222( .a(s1[21]), .b(s1[22]), .cin(s1[23]), .sum(s2[60]), .cout(c2[60]) );
FA fa223( .a(s1[25]), .b(s1[26]), .cin(s1[27]), .sum(s2[61]), .cout(c2[61]) );
FA fa224( .a(c2[52]), .b(c2[53]), .cin(c2[54]), .sum(s2[62]), .cout(c2[62]) );
FA fa225( .a(A_reg[3] & B_reg[23]), .b(A_reg[7] & B_reg[19]), .cin(A_reg[11] & B_reg[15]), .sum(s2[63]), .cout(c2[63]) );
FA fa226( .a(A_reg[19] & B_reg[7]), .b(A_reg[23] & B_reg[3]), .cin(c1[21]), .sum(s2[64]), .cout(c2[64]) );
FA fa227( .a(c1[25]), .b(c1[26]), .cin(c1[27]), .sum(s2[65]), .cout(c2[65]) );
FA fa228( .a(s1[29]), .b(s1[30]), .cin(s1[31]), .sum(s2[66]), .cout(c2[66]) );
FA fa229( .a(s1[33]), .b(s1[34]), .cin(s1[35]), .sum(s2[67]), .cout(c2[67]) );
FA fa230( .a(c2[58]), .b(c2[59]), .cin(c2[60]), .sum(s2[68]), .cout(c2[68]) );
FA fa231( .a(A_reg[3] & B_reg[24]), .b(A_reg[7] & B_reg[20]), .cin(A_reg[11] & B_reg[16]), .sum(s2[69]), .cout(c2[69]) );
FA fa232( .a(A_reg[19] & B_reg[8]), .b(A_reg[23] & B_reg[4]), .cin(A_reg[27] & B_reg[0]), .sum(s2[70]), .cout(c2[70]) );
FA fa233( .a(c1[34]), .b(c1[35]), .cin(s1[36]), .sum(s2[71]), .cout(c2[71]) );
FA fa234( .a(s1[38]), .b(s1[39]), .cin(s1[40]), .sum(s2[72]), .cout(c2[72]) );
FA fa235( .a(s1[42]), .b(s1[43]), .cin(s1[44]), .sum(s2[73]), .cout(c2[73]) );
FA fa236( .a(c2[64]), .b(c2[65]), .cin(c2[66]), .sum(s2[74]), .cout(c2[74]) );
FA fa237( .a(A_reg[5] & B_reg[23]), .b(A_reg[9] & B_reg[19]), .cin(A_reg[13] & B_reg[15]), .sum(s2[75]), .cout(c2[75]) );
FA fa238( .a(A_reg[21] & B_reg[7]), .b(A_reg[25] & B_reg[3]), .cin(s0[0]), .sum(s2[76]), .cout(c2[76]) );
FA fa239( .a(c1[43]), .b(c1[44]), .cin(s1[45]), .sum(s2[77]), .cout(c2[77]) );
FA fa240( .a(s1[47]), .b(s1[48]), .cin(s1[49]), .sum(s2[78]), .cout(c2[78]) );
FA fa241( .a(s1[51]), .b(s1[52]), .cin(s1[53]), .sum(s2[79]), .cout(c2[79]) );
FA fa242( .a(c2[70]), .b(c2[71]), .cin(c2[72]), .sum(s2[80]), .cout(c2[80]) );
FA fa243( .a(A_reg[8] & B_reg[21]), .b(A_reg[12] & B_reg[17]), .cin(A_reg[16] & B_reg[13]), .sum(s2[81]), .cout(c2[81]) );
FA fa244( .a(A_reg[24] & B_reg[5]), .b(A_reg[28] & B_reg[1]), .cin(s0[2]), .sum(s2[82]), .cout(c2[82]) );
FA fa245( .a(c1[52]), .b(c1[53]), .cin(s1[54]), .sum(s2[83]), .cout(c2[83]) );
FA fa246( .a(s1[56]), .b(s1[57]), .cin(s1[58]), .sum(s2[84]), .cout(c2[84]) );
FA fa247( .a(s1[60]), .b(s1[61]), .cin(s1[62]), .sum(s2[85]), .cout(c2[85]) );
FA fa248( .a(c2[76]), .b(c2[77]), .cin(c2[78]), .sum(s2[86]), .cout(c2[86]) );
FA fa249( .a(A_reg[11] & B_reg[19]), .b(A_reg[15] & B_reg[15]), .cin(A_reg[19] & B_reg[11]), .sum(s2[87]), .cout(c2[87]) );
FA fa250( .a(A_reg[27] & B_reg[3]), .b(c0[1]), .cin(s0[5]), .sum(s2[88]), .cout(c2[88]) );
FA fa251( .a(c1[61]), .b(c1[62]), .cin(s1[63]), .sum(s2[89]), .cout(c2[89]) );
FA fa252( .a(s1[65]), .b(s1[66]), .cin(s1[67]), .sum(s2[90]), .cout(c2[90]) );
FA fa253( .a(s1[69]), .b(s1[70]), .cin(s1[71]), .sum(s2[91]), .cout(c2[91]) );
FA fa254( .a(c2[82]), .b(c2[83]), .cin(c2[84]), .sum(s2[92]), .cout(c2[92]) );
FA fa255( .a(A_reg[14] & B_reg[17]), .b(A_reg[18] & B_reg[13]), .cin(A_reg[22] & B_reg[9]), .sum(s2[93]), .cout(c2[93]) );
FA fa256( .a(A_reg[30] & B_reg[1]), .b(c0[5]), .cin(s0[9]), .sum(s2[94]), .cout(c2[94]) );
FA fa257( .a(c1[70]), .b(c1[71]), .cin(s1[72]), .sum(s2[95]), .cout(c2[95]) );
FA fa258( .a(s1[74]), .b(s1[75]), .cin(s1[76]), .sum(s2[96]), .cout(c2[96]) );
FA fa259( .a(s1[78]), .b(s1[79]), .cin(s1[80]), .sum(s2[97]), .cout(c2[97]) );
FA fa260( .a(c2[88]), .b(c2[89]), .cin(c2[90]), .sum(s2[98]), .cout(c2[98]) );
FA fa261( .a(A_reg[15] & B_reg[17]), .b(A_reg[19] & B_reg[13]), .cin(A_reg[23] & B_reg[9]), .sum(s2[99]), .cout(c2[99]) );
FA fa262( .a(A_reg[31] & B_reg[1]), .b(c0[9]), .cin(s0[13]), .sum(s2[100]), .cout(c2[100]) );
FA fa263( .a(c1[79]), .b(c1[80]), .cin(s1[81]), .sum(s2[101]), .cout(c2[101]) );
FA fa264( .a(s1[83]), .b(s1[84]), .cin(s1[85]), .sum(s2[102]), .cout(c2[102]) );
FA fa265( .a(s1[87]), .b(s1[88]), .cin(s1[89]), .sum(s2[103]), .cout(c2[103]) );
FA fa266( .a(c2[94]), .b(c2[95]), .cin(c2[96]), .sum(s2[104]), .cout(c2[104]) );
FA fa267( .a(A_reg[14] & B_reg[19]), .b(A_reg[18] & B_reg[15]), .cin(A_reg[22] & B_reg[11]), .sum(s2[105]), .cout(c2[105]) );
FA fa268( .a(A_reg[30] & B_reg[3]), .b(c0[12]), .cin(s0[16]), .sum(s2[106]), .cout(c2[106]) );
FA fa269( .a(c1[88]), .b(c1[89]), .cin(s1[90]), .sum(s2[107]), .cout(c2[107]) );
FA fa270( .a(s1[92]), .b(s1[93]), .cin(s1[94]), .sum(s2[108]), .cout(c2[108]) );
FA fa271( .a(s1[96]), .b(s1[97]), .cin(s1[98]), .sum(s2[109]), .cout(c2[109]) );
FA fa272( .a(c2[100]), .b(c2[101]), .cin(c2[102]), .sum(s2[110]), .cout(c2[110]) );
FA fa273( .a(A_reg[12] & B_reg[22]), .b(A_reg[16] & B_reg[18]), .cin(A_reg[20] & B_reg[14]), .sum(s2[111]), .cout(c2[111]) );
FA fa274( .a(A_reg[28] & B_reg[6]), .b(c0[14]), .cin(s0[18]), .sum(s2[112]), .cout(c2[112]) );
FA fa275( .a(c1[97]), .b(c1[98]), .cin(s1[99]), .sum(s2[113]), .cout(c2[113]) );
FA fa276( .a(s1[101]), .b(s1[102]), .cin(s1[103]), .sum(s2[114]), .cout(c2[114]) );
FA fa277( .a(s1[105]), .b(s1[106]), .cin(s1[107]), .sum(s2[115]), .cout(c2[115]) );
FA fa278( .a(c2[106]), .b(c2[107]), .cin(c2[108]), .sum(s2[116]), .cout(c2[116]) );
FA fa279( .a(A_reg[10] & B_reg[25]), .b(A_reg[14] & B_reg[21]), .cin(A_reg[18] & B_reg[17]), .sum(s2[117]), .cout(c2[117]) );
FA fa280( .a(A_reg[26] & B_reg[9]), .b(A_reg[30] & B_reg[5]), .cin(s0[19]), .sum(s2[118]), .cout(c2[118]) );
FA fa281( .a(c1[106]), .b(c1[107]), .cin(s1[108]), .sum(s2[119]), .cout(c2[119]) );
FA fa282( .a(s1[110]), .b(s1[111]), .cin(s1[112]), .sum(s2[120]), .cout(c2[120]) );
FA fa283( .a(s1[114]), .b(s1[115]), .cin(s1[116]), .sum(s2[121]), .cout(c2[121]) );
FA fa284( .a(c2[112]), .b(c2[113]), .cin(c2[114]), .sum(s2[122]), .cout(c2[122]) );
FA fa285( .a(A_reg[8] & B_reg[28]), .b(A_reg[12] & B_reg[24]), .cin(A_reg[16] & B_reg[20]), .sum(s2[123]), .cout(c2[123]) );
FA fa286( .a(A_reg[24] & B_reg[12]), .b(A_reg[28] & B_reg[8]), .cin(c0[19]), .sum(s2[124]), .cout(c2[124]) );
FA fa287( .a(c1[115]), .b(c1[116]), .cin(s1[117]), .sum(s2[125]), .cout(c2[125]) );
FA fa288( .a(s1[119]), .b(s1[120]), .cin(s1[121]), .sum(s2[126]), .cout(c2[126]) );
FA fa289( .a(s1[123]), .b(s1[124]), .cin(s1[125]), .sum(s2[127]), .cout(c2[127]) );
FA fa290( .a(c2[118]), .b(c2[119]), .cin(c2[120]), .sum(s2[128]), .cout(c2[128]) );
FA fa291( .a(A_reg[9] & B_reg[28]), .b(A_reg[13] & B_reg[24]), .cin(A_reg[17] & B_reg[20]), .sum(s2[129]), .cout(c2[129]) );
FA fa292( .a(A_reg[25] & B_reg[12]), .b(A_reg[29] & B_reg[8]), .cin(c1[118]), .sum(s2[130]), .cout(c2[130]) );
FA fa293( .a(c1[123]), .b(c1[124]), .cin(c1[125]), .sum(s2[131]), .cout(c2[131]) );
FA fa294( .a(s1[127]), .b(s1[128]), .cin(s1[129]), .sum(s2[132]), .cout(c2[132]) );
FA fa295( .a(s1[131]), .b(s1[132]), .cin(s1[133]), .sum(s2[133]), .cout(c2[133]) );
FA fa296( .a(c2[124]), .b(c2[125]), .cin(c2[126]), .sum(s2[134]), .cout(c2[134]) );
FA fa297( .a(A_reg[10] & B_reg[28]), .b(A_reg[14] & B_reg[24]), .cin(A_reg[18] & B_reg[20]), .sum(s2[135]), .cout(c2[135]) );
FA fa298( .a(A_reg[26] & B_reg[12]), .b(A_reg[30] & B_reg[8]), .cin(c1[128]), .sum(s2[136]), .cout(c2[136]) );
FA fa299( .a(c1[130]), .b(c1[131]), .cin(c1[132]), .sum(s2[137]), .cout(c2[137]) );
FA fa300( .a(s1[134]), .b(s1[135]), .cin(s1[136]), .sum(s2[138]), .cout(c2[138]) );
FA fa301( .a(s1[138]), .b(s1[139]), .cin(s1[140]), .sum(s2[139]), .cout(c2[139]) );
FA fa302( .a(c2[130]), .b(c2[131]), .cin(c2[132]), .sum(s2[140]), .cout(c2[140]) );
FA fa303( .a(A_reg[11] & B_reg[28]), .b(A_reg[15] & B_reg[24]), .cin(A_reg[19] & B_reg[20]), .sum(s2[141]), .cout(c2[141]) );
FA fa304( .a(A_reg[27] & B_reg[12]), .b(A_reg[31] & B_reg[8]), .cin(c1[134]), .sum(s2[142]), .cout(c2[142]) );
FA fa305( .a(c1[136]), .b(c1[137]), .cin(c1[138]), .sum(s2[143]), .cout(c2[143]) );
FA fa306( .a(c1[140]), .b(s1[141]), .cin(s1[142]), .sum(s2[144]), .cout(c2[144]) );
FA fa307( .a(s1[144]), .b(s1[145]), .cin(s1[146]), .sum(s2[145]), .cout(c2[145]) );
FA fa308( .a(c2[136]), .b(c2[137]), .cin(c2[138]), .sum(s2[146]), .cout(c2[146]) );
FA fa309( .a(A_reg[12] & B_reg[28]), .b(A_reg[16] & B_reg[24]), .cin(A_reg[20] & B_reg[20]), .sum(s2[147]), .cout(c2[147]) );
FA fa310( .a(A_reg[28] & B_reg[12]), .b(A_reg[29] & B_reg[11]), .cin(A_reg[30] & B_reg[10]), .sum(s2[148]), .cout(c2[148]) );
FA fa311( .a(c1[141]), .b(c1[142]), .cin(c1[143]), .sum(s2[149]), .cout(c2[149]) );
FA fa312( .a(c1[145]), .b(c1[146]), .cin(s1[147]), .sum(s2[150]), .cout(c2[150]) );
FA fa313( .a(s1[149]), .b(s1[150]), .cin(s1[151]), .sum(s2[151]), .cout(c2[151]) );
FA fa314( .a(c2[142]), .b(c2[143]), .cin(c2[144]), .sum(s2[152]), .cout(c2[152]) );
FA fa315( .a(A_reg[13] & B_reg[28]), .b(A_reg[17] & B_reg[24]), .cin(A_reg[21] & B_reg[20]), .sum(s2[153]), .cout(c2[153]) );
FA fa316( .a(A_reg[26] & B_reg[15]), .b(A_reg[27] & B_reg[14]), .cin(A_reg[28] & B_reg[13]), .sum(s2[154]), .cout(c2[154]) );
FA fa317( .a(A_reg[30] & B_reg[11]), .b(A_reg[31] & B_reg[10]), .cin(c1[147]), .sum(s2[155]), .cout(c2[155]) );
FA fa318( .a(c1[149]), .b(c1[150]), .cin(c1[151]), .sum(s2[156]), .cout(c2[156]) );
FA fa319( .a(s1[153]), .b(s1[154]), .cin(s1[155]), .sum(s2[157]), .cout(c2[157]) );
FA fa320( .a(c2[148]), .b(c2[149]), .cin(c2[150]), .sum(s2[158]), .cout(c2[158]) );
FA fa321( .a(A_reg[14] & B_reg[28]), .b(A_reg[18] & B_reg[24]), .cin(A_reg[22] & B_reg[20]), .sum(s2[159]), .cout(c2[159]) );
FA fa322( .a(A_reg[24] & B_reg[18]), .b(A_reg[25] & B_reg[17]), .cin(A_reg[26] & B_reg[16]), .sum(s2[160]), .cout(c2[160]) );
FA fa323( .a(A_reg[28] & B_reg[14]), .b(A_reg[29] & B_reg[13]), .cin(A_reg[30] & B_reg[12]), .sum(s2[161]), .cout(c2[161]) );
FA fa324( .a(c1[152]), .b(c1[153]), .cin(c1[154]), .sum(s2[162]), .cout(c2[162]) );
FA fa325( .a(s1[156]), .b(s1[157]), .cin(s1[158]), .sum(s2[163]), .cout(c2[163]) );
FA fa326( .a(c2[154]), .b(c2[155]), .cin(c2[156]), .sum(s2[164]), .cout(c2[164]) );
FA fa327( .a(A_reg[15] & B_reg[28]), .b(A_reg[19] & B_reg[24]), .cin(A_reg[20] & B_reg[23]), .sum(s2[165]), .cout(c2[165]) );
FA fa328( .a(A_reg[22] & B_reg[21]), .b(A_reg[23] & B_reg[20]), .cin(A_reg[24] & B_reg[19]), .sum(s2[166]), .cout(c2[166]) );
FA fa329( .a(A_reg[26] & B_reg[17]), .b(A_reg[27] & B_reg[16]), .cin(A_reg[28] & B_reg[15]), .sum(s2[167]), .cout(c2[167]) );
FA fa330( .a(A_reg[30] & B_reg[13]), .b(A_reg[31] & B_reg[12]), .cin(c1[156]), .sum(s2[168]), .cout(c2[168]) );
FA fa331( .a(c1[158]), .b(s1[159]), .cin(s1[160]), .sum(s2[169]), .cout(c2[169]) );
FA fa332( .a(c2[160]), .b(c2[161]), .cin(c2[162]), .sum(s2[170]), .cout(c2[170]) );
FA fa333( .a(A_reg[16] & B_reg[28]), .b(A_reg[17] & B_reg[27]), .cin(A_reg[18] & B_reg[26]), .sum(s2[171]), .cout(c2[171]) );
FA fa334( .a(A_reg[20] & B_reg[24]), .b(A_reg[21] & B_reg[23]), .cin(A_reg[22] & B_reg[22]), .sum(s2[172]), .cout(c2[172]) );
FA fa335( .a(A_reg[24] & B_reg[20]), .b(A_reg[25] & B_reg[19]), .cin(A_reg[26] & B_reg[18]), .sum(s2[173]), .cout(c2[173]) );
FA fa336( .a(A_reg[28] & B_reg[16]), .b(A_reg[29] & B_reg[15]), .cin(A_reg[30] & B_reg[14]), .sum(s2[174]), .cout(c2[174]) );
FA fa337( .a(c1[159]), .b(c1[160]), .cin(s1[161]), .sum(s2[175]), .cout(c2[175]) );
FA fa338( .a(c2[166]), .b(c2[167]), .cin(c2[168]), .sum(s2[176]), .cout(c2[176]) );
FA fa339( .a(A_reg[14] & B_reg[31]), .b(A_reg[15] & B_reg[30]), .cin(A_reg[16] & B_reg[29]), .sum(s2[177]), .cout(c2[177]) );
FA fa340( .a(A_reg[18] & B_reg[27]), .b(A_reg[19] & B_reg[26]), .cin(A_reg[20] & B_reg[25]), .sum(s2[178]), .cout(c2[178]) );
FA fa341( .a(A_reg[22] & B_reg[23]), .b(A_reg[23] & B_reg[22]), .cin(A_reg[24] & B_reg[21]), .sum(s2[179]), .cout(c2[179]) );
FA fa342( .a(A_reg[26] & B_reg[19]), .b(A_reg[27] & B_reg[18]), .cin(A_reg[28] & B_reg[17]), .sum(s2[180]), .cout(c2[180]) );
FA fa343( .a(A_reg[30] & B_reg[15]), .b(A_reg[31] & B_reg[14]), .cin(c1[161]), .sum(s2[181]), .cout(c2[181]) );
FA fa344( .a(c2[172]), .b(c2[173]), .cin(c2[174]), .sum(s2[182]), .cout(c2[182]) );
FA fa345( .a(A_reg[15] & B_reg[31]), .b(A_reg[16] & B_reg[30]), .cin(A_reg[17] & B_reg[29]), .sum(s2[183]), .cout(c2[183]) );
FA fa346( .a(A_reg[19] & B_reg[27]), .b(A_reg[20] & B_reg[26]), .cin(A_reg[21] & B_reg[25]), .sum(s2[184]), .cout(c2[184]) );
FA fa347( .a(A_reg[23] & B_reg[23]), .b(A_reg[24] & B_reg[22]), .cin(A_reg[25] & B_reg[21]), .sum(s2[185]), .cout(c2[185]) );
FA fa348( .a(A_reg[27] & B_reg[19]), .b(A_reg[28] & B_reg[18]), .cin(A_reg[29] & B_reg[17]), .sum(s2[186]), .cout(c2[186]) );
FA fa349( .a(A_reg[31] & B_reg[15]), .b(c2[177]), .cin(c2[178]), .sum(s2[187]), .cout(c2[187]) );
FA fa350( .a(A_reg[16] & B_reg[31]), .b(A_reg[17] & B_reg[30]), .cin(A_reg[18] & B_reg[29]), .sum(s2[188]), .cout(c2[188]) );
FA fa351( .a(A_reg[20] & B_reg[27]), .b(A_reg[21] & B_reg[26]), .cin(A_reg[22] & B_reg[25]), .sum(s2[189]), .cout(c2[189]) );
FA fa352( .a(A_reg[24] & B_reg[23]), .b(A_reg[25] & B_reg[22]), .cin(A_reg[26] & B_reg[21]), .sum(s2[190]), .cout(c2[190]) );
FA fa353( .a(A_reg[28] & B_reg[19]), .b(A_reg[29] & B_reg[18]), .cin(A_reg[30] & B_reg[17]), .sum(s2[191]), .cout(c2[191]) );
FA fa354( .a(A_reg[17] & B_reg[31]), .b(A_reg[18] & B_reg[30]), .cin(A_reg[19] & B_reg[29]), .sum(s2[192]), .cout(c2[192]) );
FA fa355( .a(A_reg[21] & B_reg[27]), .b(A_reg[22] & B_reg[26]), .cin(A_reg[23] & B_reg[25]), .sum(s2[193]), .cout(c2[193]) );
FA fa356( .a(A_reg[25] & B_reg[23]), .b(A_reg[26] & B_reg[22]), .cin(A_reg[27] & B_reg[21]), .sum(s2[194]), .cout(c2[194]) );
FA fa357( .a(A_reg[18] & B_reg[31]), .b(A_reg[19] & B_reg[30]), .cin(A_reg[20] & B_reg[29]), .sum(s2[195]), .cout(c2[195]) );
FA fa358( .a(A_reg[22] & B_reg[27]), .b(A_reg[23] & B_reg[26]), .cin(A_reg[24] & B_reg[25]), .sum(s2[196]), .cout(c2[196]) );
FA fa359( .a(A_reg[19] & B_reg[31]), .b(A_reg[20] & B_reg[30]), .cin(A_reg[21] & B_reg[29]), .sum(s2[197]), .cout(c2[197]) );
//stage 3 reduction
HA ha20( .a(A_reg[0] & B_reg[9]), .b(A_reg[1] & B_reg[8]), .sum(s3[0]), .cout(c3[0]) );
FA fa360( .a(A_reg[0] & B_reg[10]), .b(A_reg[1] & B_reg[9]), .cin(A_reg[2] & B_reg[8]), .sum(s3[1]), .cout(c3[1]) );
HA ha21( .a(A_reg[4] & B_reg[6]), .b(A_reg[5] & B_reg[5]), .sum(s3[2]), .cout(c3[2]) );
FA fa361( .a(A_reg[0] & B_reg[11]), .b(A_reg[1] & B_reg[10]), .cin(A_reg[2] & B_reg[9]), .sum(s3[3]), .cout(c3[3]) );
FA fa362( .a(A_reg[4] & B_reg[7]), .b(A_reg[5] & B_reg[6]), .cin(A_reg[6] & B_reg[5]), .sum(s3[4]), .cout(c3[4]) );
HA ha22( .a(A_reg[8] & B_reg[3]), .b(A_reg[9] & B_reg[2]), .sum(s3[5]), .cout(c3[5]) );
FA fa363( .a(A_reg[0] & B_reg[12]), .b(A_reg[1] & B_reg[11]), .cin(A_reg[2] & B_reg[10]), .sum(s3[6]), .cout(c3[6]) );
FA fa364( .a(A_reg[4] & B_reg[8]), .b(A_reg[5] & B_reg[7]), .cin(A_reg[6] & B_reg[6]), .sum(s3[7]), .cout(c3[7]) );
FA fa365( .a(A_reg[8] & B_reg[4]), .b(A_reg[9] & B_reg[3]), .cin(A_reg[10] & B_reg[2]), .sum(s3[8]), .cout(c3[8]) );
HA ha23( .a(A_reg[12] & B_reg[0]), .b(c3[3]), .sum(s3[9]), .cout(c3[9]) );
FA fa366( .a(A_reg[2] & B_reg[11]), .b(A_reg[3] & B_reg[10]), .cin(A_reg[4] & B_reg[9]), .sum(s3[10]), .cout(c3[10]) );
FA fa367( .a(A_reg[6] & B_reg[7]), .b(A_reg[7] & B_reg[6]), .cin(A_reg[8] & B_reg[5]), .sum(s3[11]), .cout(c3[11]) );
FA fa368( .a(A_reg[10] & B_reg[3]), .b(A_reg[11] & B_reg[2]), .cin(A_reg[12] & B_reg[1]), .sum(s3[12]), .cout(c3[12]) );
FA fa369( .a(s2[0]), .b(c3[6]), .cin(c3[7]), .sum(s3[13]), .cout(c3[13]) );
FA fa370( .a(A_reg[3] & B_reg[11]), .b(A_reg[6] & B_reg[8]), .cin(A_reg[7] & B_reg[7]), .sum(s3[14]), .cout(c3[14]) );
FA fa371( .a(A_reg[9] & B_reg[5]), .b(A_reg[10] & B_reg[4]), .cin(A_reg[11] & B_reg[3]), .sum(s3[15]), .cout(c3[15]) );
FA fa372( .a(A_reg[13] & B_reg[1]), .b(A_reg[14] & B_reg[0]), .cin(c2[0]), .sum(s3[16]), .cout(c3[16]) );
FA fa373( .a(s2[2]), .b(c3[10]), .cin(c3[11]), .sum(s3[17]), .cout(c3[17]) );
FA fa374( .a(A_reg[3] & B_reg[12]), .b(A_reg[7] & B_reg[8]), .cin(A_reg[10] & B_reg[5]), .sum(s3[18]), .cout(c3[18]) );
FA fa375( .a(A_reg[12] & B_reg[3]), .b(A_reg[13] & B_reg[2]), .cin(A_reg[14] & B_reg[1]), .sum(s3[19]), .cout(c3[19]) );
FA fa376( .a(c2[1]), .b(c2[2]), .cin(s2[3]), .sum(s3[20]), .cout(c3[20]) );
FA fa377( .a(s2[5]), .b(c3[14]), .cin(c3[15]), .sum(s3[21]), .cout(c3[21]) );
FA fa378( .a(A_reg[3] & B_reg[13]), .b(A_reg[7] & B_reg[9]), .cin(A_reg[11] & B_reg[5]), .sum(s3[22]), .cout(c3[22]) );
FA fa379( .a(A_reg[15] & B_reg[1]), .b(A_reg[16] & B_reg[0]), .cin(c2[3]), .sum(s3[23]), .cout(c3[23]) );
FA fa380( .a(c2[5]), .b(s2[6]), .cin(s2[7]), .sum(s3[24]), .cout(c3[24]) );
FA fa381( .a(s2[9]), .b(c3[18]), .cin(c3[19]), .sum(s3[25]), .cout(c3[25]) );
FA fa382( .a(A_reg[3] & B_reg[14]), .b(A_reg[7] & B_reg[10]), .cin(A_reg[11] & B_reg[6]), .sum(s3[26]), .cout(c3[26]) );
FA fa383( .a(c2[6]), .b(c2[7]), .cin(c2[8]), .sum(s3[27]), .cout(c3[27]) );
FA fa384( .a(s2[10]), .b(s2[11]), .cin(s2[12]), .sum(s3[28]), .cout(c3[28]) );
FA fa385( .a(s2[14]), .b(c3[22]), .cin(c3[23]), .sum(s3[29]), .cout(c3[29]) );
FA fa386( .a(A_reg[3] & B_reg[15]), .b(A_reg[7] & B_reg[11]), .cin(A_reg[11] & B_reg[7]), .sum(s3[30]), .cout(c3[30]) );
FA fa387( .a(c2[10]), .b(c2[13]), .cin(c2[14]), .sum(s3[31]), .cout(c3[31]) );
FA fa388( .a(s2[16]), .b(s2[17]), .cin(s2[18]), .sum(s3[32]), .cout(c3[32]) );
FA fa389( .a(s2[20]), .b(c3[26]), .cin(c3[27]), .sum(s3[33]), .cout(c3[33]) );
FA fa390( .a(A_reg[5] & B_reg[14]), .b(A_reg[9] & B_reg[10]), .cin(A_reg[13] & B_reg[6]), .sum(s3[34]), .cout(c3[34]) );
FA fa391( .a(c2[15]), .b(c2[19]), .cin(c2[20]), .sum(s3[35]), .cout(c3[35]) );
FA fa392( .a(s2[22]), .b(s2[23]), .cin(s2[24]), .sum(s3[36]), .cout(c3[36]) );
FA fa393( .a(s2[26]), .b(c3[30]), .cin(c3[31]), .sum(s3[37]), .cout(c3[37]) );
FA fa394( .a(A_reg[8] & B_reg[12]), .b(A_reg[12] & B_reg[8]), .cin(A_reg[16] & B_reg[4]), .sum(s3[38]), .cout(c3[38]) );
FA fa395( .a(c2[21]), .b(c2[25]), .cin(c2[26]), .sum(s3[39]), .cout(c3[39]) );
FA fa396( .a(s2[28]), .b(s2[29]), .cin(s2[30]), .sum(s3[40]), .cout(c3[40]) );
FA fa397( .a(s2[32]), .b(c3[34]), .cin(c3[35]), .sum(s3[41]), .cout(c3[41]) );
FA fa398( .a(A_reg[11] & B_reg[10]), .b(A_reg[15] & B_reg[6]), .cin(A_reg[19] & B_reg[2]), .sum(s3[42]), .cout(c3[42]) );
FA fa399( .a(c2[27]), .b(c2[31]), .cin(c2[32]), .sum(s3[43]), .cout(c3[43]) );
FA fa400( .a(s2[34]), .b(s2[35]), .cin(s2[36]), .sum(s3[44]), .cout(c3[44]) );
FA fa401( .a(s2[38]), .b(c3[38]), .cin(c3[39]), .sum(s3[45]), .cout(c3[45]) );
FA fa402( .a(A_reg[14] & B_reg[8]), .b(A_reg[18] & B_reg[4]), .cin(A_reg[22] & B_reg[0]), .sum(s3[46]), .cout(c3[46]) );
FA fa403( .a(c2[33]), .b(c2[37]), .cin(c2[38]), .sum(s3[47]), .cout(c3[47]) );
FA fa404( .a(s2[40]), .b(s2[41]), .cin(s2[42]), .sum(s3[48]), .cout(c3[48]) );
FA fa405( .a(s2[44]), .b(c3[42]), .cin(c3[43]), .sum(s3[49]), .cout(c3[49]) );
FA fa406( .a(A_reg[15] & B_reg[8]), .b(A_reg[21] & B_reg[2]), .cin(c1[7]), .sum(s3[50]), .cout(c3[50]) );
FA fa407( .a(c2[39]), .b(c2[43]), .cin(c2[44]), .sum(s3[51]), .cout(c3[51]) );
FA fa408( .a(s2[46]), .b(s2[47]), .cin(s2[48]), .sum(s3[52]), .cout(c3[52]) );
FA fa409( .a(s2[50]), .b(c3[46]), .cin(c3[47]), .sum(s3[53]), .cout(c3[53]) );
FA fa410( .a(A_reg[15] & B_reg[9]), .b(A_reg[24] & B_reg[0]), .cin(c1[13]), .sum(s3[54]), .cout(c3[54]) );
FA fa411( .a(c2[45]), .b(c2[49]), .cin(c2[50]), .sum(s3[55]), .cout(c3[55]) );
FA fa412( .a(s2[52]), .b(s2[53]), .cin(s2[54]), .sum(s3[56]), .cout(c3[56]) );
FA fa413( .a(s2[56]), .b(c3[50]), .cin(c3[51]), .sum(s3[57]), .cout(c3[57]) );
FA fa414( .a(A_reg[15] & B_reg[10]), .b(c1[16]), .cin(c1[20]), .sum(s3[58]), .cout(c3[58]) );
FA fa415( .a(c2[51]), .b(c2[55]), .cin(c2[56]), .sum(s3[59]), .cout(c3[59]) );
FA fa416( .a(s2[58]), .b(s2[59]), .cin(s2[60]), .sum(s3[60]), .cout(c3[60]) );
FA fa417( .a(s2[62]), .b(c3[54]), .cin(c3[55]), .sum(s3[61]), .cout(c3[61]) );
FA fa418( .a(A_reg[15] & B_reg[11]), .b(c1[24]), .cin(s1[28]), .sum(s3[62]), .cout(c3[62]) );
FA fa419( .a(c2[57]), .b(c2[61]), .cin(c2[62]), .sum(s3[63]), .cout(c3[63]) );
FA fa420( .a(s2[64]), .b(s2[65]), .cin(s2[66]), .sum(s3[64]), .cout(c3[64]) );
FA fa421( .a(s2[68]), .b(c3[58]), .cin(c3[59]), .sum(s3[65]), .cout(c3[65]) );
FA fa422( .a(A_reg[15] & B_reg[12]), .b(c1[31]), .cin(s1[37]), .sum(s3[66]), .cout(c3[66]) );
FA fa423( .a(c2[63]), .b(c2[67]), .cin(c2[68]), .sum(s3[67]), .cout(c3[67]) );
FA fa424( .a(s2[70]), .b(s2[71]), .cin(s2[72]), .sum(s3[68]), .cout(c3[68]) );
FA fa425( .a(s2[74]), .b(c3[62]), .cin(c3[63]), .sum(s3[69]), .cout(c3[69]) );
FA fa426( .a(A_reg[17] & B_reg[11]), .b(c1[39]), .cin(s1[46]), .sum(s3[70]), .cout(c3[70]) );
FA fa427( .a(c2[69]), .b(c2[73]), .cin(c2[74]), .sum(s3[71]), .cout(c3[71]) );
FA fa428( .a(s2[76]), .b(s2[77]), .cin(s2[78]), .sum(s3[72]), .cout(c3[72]) );
FA fa429( .a(s2[80]), .b(c3[66]), .cin(c3[67]), .sum(s3[73]), .cout(c3[73]) );
FA fa430( .a(A_reg[20] & B_reg[9]), .b(c1[48]), .cin(s1[55]), .sum(s3[74]), .cout(c3[74]) );
FA fa431( .a(c2[75]), .b(c2[79]), .cin(c2[80]), .sum(s3[75]), .cout(c3[75]) );
FA fa432( .a(s2[82]), .b(s2[83]), .cin(s2[84]), .sum(s3[76]), .cout(c3[76]) );
FA fa433( .a(s2[86]), .b(c3[70]), .cin(c3[71]), .sum(s3[77]), .cout(c3[77]) );
FA fa434( .a(A_reg[23] & B_reg[7]), .b(c1[57]), .cin(s1[64]), .sum(s3[78]), .cout(c3[78]) );
FA fa435( .a(c2[81]), .b(c2[85]), .cin(c2[86]), .sum(s3[79]), .cout(c3[79]) );
FA fa436( .a(s2[88]), .b(s2[89]), .cin(s2[90]), .sum(s3[80]), .cout(c3[80]) );
FA fa437( .a(s2[92]), .b(c3[74]), .cin(c3[75]), .sum(s3[81]), .cout(c3[81]) );
FA fa438( .a(A_reg[26] & B_reg[5]), .b(c1[66]), .cin(s1[73]), .sum(s3[82]), .cout(c3[82]) );
FA fa439( .a(c2[87]), .b(c2[91]), .cin(c2[92]), .sum(s3[83]), .cout(c3[83]) );
FA fa440( .a(s2[94]), .b(s2[95]), .cin(s2[96]), .sum(s3[84]), .cout(c3[84]) );
FA fa441( .a(s2[98]), .b(c3[78]), .cin(c3[79]), .sum(s3[85]), .cout(c3[85]) );
FA fa442( .a(A_reg[27] & B_reg[5]), .b(c1[75]), .cin(s1[82]), .sum(s3[86]), .cout(c3[86]) );
FA fa443( .a(c2[93]), .b(c2[97]), .cin(c2[98]), .sum(s3[87]), .cout(c3[87]) );
FA fa444( .a(s2[100]), .b(s2[101]), .cin(s2[102]), .sum(s3[88]), .cout(c3[88]) );
FA fa445( .a(s2[104]), .b(c3[82]), .cin(c3[83]), .sum(s3[89]), .cout(c3[89]) );
FA fa446( .a(A_reg[26] & B_reg[7]), .b(c1[84]), .cin(s1[91]), .sum(s3[90]), .cout(c3[90]) );
FA fa447( .a(c2[99]), .b(c2[103]), .cin(c2[104]), .sum(s3[91]), .cout(c3[91]) );
FA fa448( .a(s2[106]), .b(s2[107]), .cin(s2[108]), .sum(s3[92]), .cout(c3[92]) );
FA fa449( .a(s2[110]), .b(c3[86]), .cin(c3[87]), .sum(s3[93]), .cout(c3[93]) );
FA fa450( .a(A_reg[24] & B_reg[10]), .b(c1[93]), .cin(s1[100]), .sum(s3[94]), .cout(c3[94]) );
FA fa451( .a(c2[105]), .b(c2[109]), .cin(c2[110]), .sum(s3[95]), .cout(c3[95]) );
FA fa452( .a(s2[112]), .b(s2[113]), .cin(s2[114]), .sum(s3[96]), .cout(c3[96]) );
FA fa453( .a(s2[116]), .b(c3[90]), .cin(c3[91]), .sum(s3[97]), .cout(c3[97]) );
FA fa454( .a(A_reg[22] & B_reg[13]), .b(c1[102]), .cin(s1[109]), .sum(s3[98]), .cout(c3[98]) );
FA fa455( .a(c2[111]), .b(c2[115]), .cin(c2[116]), .sum(s3[99]), .cout(c3[99]) );
FA fa456( .a(s2[118]), .b(s2[119]), .cin(s2[120]), .sum(s3[100]), .cout(c3[100]) );
FA fa457( .a(s2[122]), .b(c3[94]), .cin(c3[95]), .sum(s3[101]), .cout(c3[101]) );
FA fa458( .a(A_reg[20] & B_reg[16]), .b(c1[111]), .cin(s1[118]), .sum(s3[102]), .cout(c3[102]) );
FA fa459( .a(c2[117]), .b(c2[121]), .cin(c2[122]), .sum(s3[103]), .cout(c3[103]) );
FA fa460( .a(s2[124]), .b(s2[125]), .cin(s2[126]), .sum(s3[104]), .cout(c3[104]) );
FA fa461( .a(s2[128]), .b(c3[98]), .cin(c3[99]), .sum(s3[105]), .cout(c3[105]) );
FA fa462( .a(A_reg[21] & B_reg[16]), .b(c1[122]), .cin(s1[126]), .sum(s3[106]), .cout(c3[106]) );
FA fa463( .a(c2[123]), .b(c2[127]), .cin(c2[128]), .sum(s3[107]), .cout(c3[107]) );
FA fa464( .a(s2[130]), .b(s2[131]), .cin(s2[132]), .sum(s3[108]), .cout(c3[108]) );
FA fa465( .a(s2[134]), .b(c3[102]), .cin(c3[103]), .sum(s3[109]), .cout(c3[109]) );
FA fa466( .a(A_reg[22] & B_reg[16]), .b(c1[129]), .cin(c1[133]), .sum(s3[110]), .cout(c3[110]) );
FA fa467( .a(c2[129]), .b(c2[133]), .cin(c2[134]), .sum(s3[111]), .cout(c3[111]) );
FA fa468( .a(s2[136]), .b(s2[137]), .cin(s2[138]), .sum(s3[112]), .cout(c3[112]) );
FA fa469( .a(s2[140]), .b(c3[106]), .cin(c3[107]), .sum(s3[113]), .cout(c3[113]) );
FA fa470( .a(A_reg[23] & B_reg[16]), .b(c1[135]), .cin(c1[139]), .sum(s3[114]), .cout(c3[114]) );
FA fa471( .a(c2[135]), .b(c2[139]), .cin(c2[140]), .sum(s3[115]), .cout(c3[115]) );
FA fa472( .a(s2[142]), .b(s2[143]), .cin(s2[144]), .sum(s3[116]), .cout(c3[116]) );
FA fa473( .a(s2[146]), .b(c3[110]), .cin(c3[111]), .sum(s3[117]), .cout(c3[117]) );
FA fa474( .a(A_reg[24] & B_reg[16]), .b(A_reg[31] & B_reg[9]), .cin(c1[144]), .sum(s3[118]), .cout(c3[118]) );
FA fa475( .a(c2[141]), .b(c2[145]), .cin(c2[146]), .sum(s3[119]), .cout(c3[119]) );
FA fa476( .a(s2[148]), .b(s2[149]), .cin(s2[150]), .sum(s3[120]), .cout(c3[120]) );
FA fa477( .a(s2[152]), .b(c3[114]), .cin(c3[115]), .sum(s3[121]), .cout(c3[121]) );
FA fa478( .a(A_reg[25] & B_reg[16]), .b(A_reg[29] & B_reg[12]), .cin(c1[148]), .sum(s3[122]), .cout(c3[122]) );
FA fa479( .a(c2[147]), .b(c2[151]), .cin(c2[152]), .sum(s3[123]), .cout(c3[123]) );
FA fa480( .a(s2[154]), .b(s2[155]), .cin(s2[156]), .sum(s3[124]), .cout(c3[124]) );
FA fa481( .a(s2[158]), .b(c3[118]), .cin(c3[119]), .sum(s3[125]), .cout(c3[125]) );
FA fa482( .a(A_reg[23] & B_reg[19]), .b(A_reg[27] & B_reg[15]), .cin(A_reg[31] & B_reg[11]), .sum(s3[126]), .cout(c3[126]) );
FA fa483( .a(c2[153]), .b(c2[157]), .cin(c2[158]), .sum(s3[127]), .cout(c3[127]) );
FA fa484( .a(s2[160]), .b(s2[161]), .cin(s2[162]), .sum(s3[128]), .cout(c3[128]) );
FA fa485( .a(s2[164]), .b(c3[122]), .cin(c3[123]), .sum(s3[129]), .cout(c3[129]) );
FA fa486( .a(A_reg[21] & B_reg[22]), .b(A_reg[25] & B_reg[18]), .cin(A_reg[29] & B_reg[14]), .sum(s3[130]), .cout(c3[130]) );
FA fa487( .a(c2[159]), .b(c2[163]), .cin(c2[164]), .sum(s3[131]), .cout(c3[131]) );
FA fa488( .a(s2[166]), .b(s2[167]), .cin(s2[168]), .sum(s3[132]), .cout(c3[132]) );
FA fa489( .a(s2[170]), .b(c3[126]), .cin(c3[127]), .sum(s3[133]), .cout(c3[133]) );
FA fa490( .a(A_reg[19] & B_reg[25]), .b(A_reg[23] & B_reg[21]), .cin(A_reg[27] & B_reg[17]), .sum(s3[134]), .cout(c3[134]) );
FA fa491( .a(c2[165]), .b(c2[169]), .cin(c2[170]), .sum(s3[135]), .cout(c3[135]) );
FA fa492( .a(s2[172]), .b(s2[173]), .cin(s2[174]), .sum(s3[136]), .cout(c3[136]) );
FA fa493( .a(s2[176]), .b(c3[130]), .cin(c3[131]), .sum(s3[137]), .cout(c3[137]) );
FA fa494( .a(A_reg[17] & B_reg[28]), .b(A_reg[21] & B_reg[24]), .cin(A_reg[25] & B_reg[20]), .sum(s3[138]), .cout(c3[138]) );
FA fa495( .a(c2[171]), .b(c2[175]), .cin(c2[176]), .sum(s3[139]), .cout(c3[139]) );
FA fa496( .a(s2[178]), .b(s2[179]), .cin(s2[180]), .sum(s3[140]), .cout(c3[140]) );
FA fa497( .a(s2[182]), .b(c3[134]), .cin(c3[135]), .sum(s3[141]), .cout(c3[141]) );
FA fa498( .a(A_reg[18] & B_reg[28]), .b(A_reg[22] & B_reg[24]), .cin(A_reg[26] & B_reg[20]), .sum(s3[142]), .cout(c3[142]) );
FA fa499( .a(c2[179]), .b(c2[180]), .cin(c2[181]), .sum(s3[143]), .cout(c3[143]) );
FA fa500( .a(s2[183]), .b(s2[184]), .cin(s2[185]), .sum(s3[144]), .cout(c3[144]) );
FA fa501( .a(s2[187]), .b(c3[138]), .cin(c3[139]), .sum(s3[145]), .cout(c3[145]) );
FA fa502( .a(A_reg[19] & B_reg[28]), .b(A_reg[23] & B_reg[24]), .cin(A_reg[27] & B_reg[20]), .sum(s3[146]), .cout(c3[146]) );
FA fa503( .a(c2[183]), .b(c2[184]), .cin(c2[185]), .sum(s3[147]), .cout(c3[147]) );
FA fa504( .a(c2[187]), .b(s2[188]), .cin(s2[189]), .sum(s3[148]), .cout(c3[148]) );
FA fa505( .a(s2[191]), .b(c3[142]), .cin(c3[143]), .sum(s3[149]), .cout(c3[149]) );
FA fa506( .a(A_reg[20] & B_reg[28]), .b(A_reg[24] & B_reg[24]), .cin(A_reg[28] & B_reg[20]), .sum(s3[150]), .cout(c3[150]) );
FA fa507( .a(A_reg[30] & B_reg[18]), .b(A_reg[31] & B_reg[17]), .cin(c2[188]), .sum(s3[151]), .cout(c3[151]) );
FA fa508( .a(c2[190]), .b(c2[191]), .cin(s2[192]), .sum(s3[152]), .cout(c3[152]) );
FA fa509( .a(s2[194]), .b(c3[146]), .cin(c3[147]), .sum(s3[153]), .cout(c3[153]) );
FA fa510( .a(A_reg[21] & B_reg[28]), .b(A_reg[25] & B_reg[24]), .cin(A_reg[26] & B_reg[23]), .sum(s3[154]), .cout(c3[154]) );
FA fa511( .a(A_reg[28] & B_reg[21]), .b(A_reg[29] & B_reg[20]), .cin(A_reg[30] & B_reg[19]), .sum(s3[155]), .cout(c3[155]) );
FA fa512( .a(c2[192]), .b(c2[193]), .cin(c2[194]), .sum(s3[156]), .cout(c3[156]) );
FA fa513( .a(s2[196]), .b(c3[150]), .cin(c3[151]), .sum(s3[157]), .cout(c3[157]) );
FA fa514( .a(A_reg[22] & B_reg[28]), .b(A_reg[23] & B_reg[27]), .cin(A_reg[24] & B_reg[26]), .sum(s3[158]), .cout(c3[158]) );
FA fa515( .a(A_reg[26] & B_reg[24]), .b(A_reg[27] & B_reg[23]), .cin(A_reg[28] & B_reg[22]), .sum(s3[159]), .cout(c3[159]) );
FA fa516( .a(A_reg[30] & B_reg[20]), .b(A_reg[31] & B_reg[19]), .cin(c2[195]), .sum(s3[160]), .cout(c3[160]) );
FA fa517( .a(s2[197]), .b(c3[154]), .cin(c3[155]), .sum(s3[161]), .cout(c3[161]) );
FA fa518( .a(A_reg[20] & B_reg[31]), .b(A_reg[21] & B_reg[30]), .cin(A_reg[22] & B_reg[29]), .sum(s3[162]), .cout(c3[162]) );
FA fa519( .a(A_reg[24] & B_reg[27]), .b(A_reg[25] & B_reg[26]), .cin(A_reg[26] & B_reg[25]), .sum(s3[163]), .cout(c3[163]) );
FA fa520( .a(A_reg[28] & B_reg[23]), .b(A_reg[29] & B_reg[22]), .cin(A_reg[30] & B_reg[21]), .sum(s3[164]), .cout(c3[164]) );
FA fa521( .a(c2[197]), .b(c3[158]), .cin(c3[159]), .sum(s3[165]), .cout(c3[165]) );
FA fa522( .a(A_reg[21] & B_reg[31]), .b(A_reg[22] & B_reg[30]), .cin(A_reg[23] & B_reg[29]), .sum(s3[166]), .cout(c3[166]) );
FA fa523( .a(A_reg[25] & B_reg[27]), .b(A_reg[26] & B_reg[26]), .cin(A_reg[27] & B_reg[25]), .sum(s3[167]), .cout(c3[167]) );
FA fa524( .a(A_reg[29] & B_reg[23]), .b(A_reg[30] & B_reg[22]), .cin(A_reg[31] & B_reg[21]), .sum(s3[168]), .cout(c3[168]) );
FA fa525( .a(A_reg[22] & B_reg[31]), .b(A_reg[23] & B_reg[30]), .cin(A_reg[24] & B_reg[29]), .sum(s3[169]), .cout(c3[169]) );
FA fa526( .a(A_reg[26] & B_reg[27]), .b(A_reg[27] & B_reg[26]), .cin(A_reg[28] & B_reg[25]), .sum(s3[170]), .cout(c3[170]) );
FA fa527( .a(A_reg[23] & B_reg[31]), .b(A_reg[24] & B_reg[30]), .cin(A_reg[25] & B_reg[29]), .sum(s3[171]), .cout(c3[171]) );
//stage 4 reduction
HA ha24( .a(A_reg[0] & B_reg[6]), .b(A_reg[1] & B_reg[5]), .sum(s4[0]), .cout(c4[0]) );
FA fa528( .a(A_reg[0] & B_reg[7]), .b(A_reg[1] & B_reg[6]), .cin(A_reg[2] & B_reg[5]), .sum(s4[1]), .cout(c4[1]) );
HA ha25( .a(A_reg[4] & B_reg[3]), .b(A_reg[5] & B_reg[2]), .sum(s4[2]), .cout(c4[2]) );
FA fa529( .a(A_reg[0] & B_reg[8]), .b(A_reg[1] & B_reg[7]), .cin(A_reg[2] & B_reg[6]), .sum(s4[3]), .cout(c4[3]) );
FA fa530( .a(A_reg[4] & B_reg[4]), .b(A_reg[5] & B_reg[3]), .cin(A_reg[6] & B_reg[2]), .sum(s4[4]), .cout(c4[4]) );
HA ha26( .a(A_reg[8] & B_reg[0]), .b(c4[1]), .sum(s4[5]), .cout(c4[5]) );
FA fa531( .a(A_reg[2] & B_reg[7]), .b(A_reg[3] & B_reg[6]), .cin(A_reg[4] & B_reg[5]), .sum(s4[6]), .cout(c4[6]) );
FA fa532( .a(A_reg[6] & B_reg[3]), .b(A_reg[7] & B_reg[2]), .cin(A_reg[8] & B_reg[1]), .sum(s4[7]), .cout(c4[7]) );
FA fa533( .a(s3[0]), .b(c4[3]), .cin(c4[4]), .sum(s4[8]), .cout(c4[8]) );
FA fa534( .a(A_reg[3] & B_reg[7]), .b(A_reg[6] & B_reg[4]), .cin(A_reg[7] & B_reg[3]), .sum(s4[9]), .cout(c4[9]) );
FA fa535( .a(A_reg[9] & B_reg[1]), .b(A_reg[10] & B_reg[0]), .cin(c3[0]), .sum(s4[10]), .cout(c4[10]) );
FA fa536( .a(s3[2]), .b(c4[6]), .cin(c4[7]), .sum(s4[11]), .cout(c4[11]) );
FA fa537( .a(A_reg[3] & B_reg[8]), .b(A_reg[7] & B_reg[4]), .cin(A_reg[10] & B_reg[1]), .sum(s4[12]), .cout(c4[12]) );
FA fa538( .a(c3[1]), .b(c3[2]), .cin(s3[3]), .sum(s4[13]), .cout(c4[13]) );
FA fa539( .a(s3[5]), .b(c4[9]), .cin(c4[10]), .sum(s4[14]), .cout(c4[14]) );
FA fa540( .a(A_reg[3] & B_reg[9]), .b(A_reg[7] & B_reg[5]), .cin(A_reg[11] & B_reg[1]), .sum(s4[15]), .cout(c4[15]) );
FA fa541( .a(c3[5]), .b(s3[6]), .cin(s3[7]), .sum(s4[16]), .cout(c4[16]) );
FA fa542( .a(s3[9]), .b(c4[12]), .cin(c4[13]), .sum(s4[17]), .cout(c4[17]) );
FA fa543( .a(A_reg[5] & B_reg[8]), .b(A_reg[9] & B_reg[4]), .cin(A_reg[13] & B_reg[0]), .sum(s4[18]), .cout(c4[18]) );
FA fa544( .a(c3[9]), .b(s3[10]), .cin(s3[11]), .sum(s4[19]), .cout(c4[19]) );
FA fa545( .a(s3[13]), .b(c4[15]), .cin(c4[16]), .sum(s4[20]), .cout(c4[20]) );
FA fa546( .a(A_reg[8] & B_reg[6]), .b(A_reg[12] & B_reg[2]), .cin(s2[1]), .sum(s4[21]), .cout(c4[21]) );
FA fa547( .a(c3[13]), .b(s3[14]), .cin(s3[15]), .sum(s4[22]), .cout(c4[22]) );
FA fa548( .a(s3[17]), .b(c4[18]), .cin(c4[19]), .sum(s4[23]), .cout(c4[23]) );
FA fa549( .a(A_reg[11] & B_reg[4]), .b(A_reg[15] & B_reg[0]), .cin(s2[4]), .sum(s4[24]), .cout(c4[24]) );
FA fa550( .a(c3[17]), .b(s3[18]), .cin(s3[19]), .sum(s4[25]), .cout(c4[25]) );
FA fa551( .a(s3[21]), .b(c4[21]), .cin(c4[22]), .sum(s4[26]), .cout(c4[26]) );
FA fa552( .a(A_reg[14] & B_reg[2]), .b(c2[4]), .cin(s2[8]), .sum(s4[27]), .cout(c4[27]) );
FA fa553( .a(c3[21]), .b(s3[22]), .cin(s3[23]), .sum(s4[28]), .cout(c4[28]) );
FA fa554( .a(s3[25]), .b(c4[24]), .cin(c4[25]), .sum(s4[29]), .cout(c4[29]) );
FA fa555( .a(A_reg[15] & B_reg[2]), .b(c2[9]), .cin(s2[13]), .sum(s4[30]), .cout(c4[30]) );
FA fa556( .a(c3[25]), .b(s3[26]), .cin(s3[27]), .sum(s4[31]), .cout(c4[31]) );
FA fa557( .a(s3[29]), .b(c4[27]), .cin(c4[28]), .sum(s4[32]), .cout(c4[32]) );
FA fa558( .a(A_reg[15] & B_reg[3]), .b(s2[15]), .cin(s2[19]), .sum(s4[33]), .cout(c4[33]) );
FA fa559( .a(c3[29]), .b(s3[30]), .cin(s3[31]), .sum(s4[34]), .cout(c4[34]) );
FA fa560( .a(s3[33]), .b(c4[30]), .cin(c4[31]), .sum(s4[35]), .cout(c4[35]) );
FA fa561( .a(A_reg[17] & B_reg[2]), .b(s2[21]), .cin(s2[25]), .sum(s4[36]), .cout(c4[36]) );
FA fa562( .a(c3[33]), .b(s3[34]), .cin(s3[35]), .sum(s4[37]), .cout(c4[37]) );
FA fa563( .a(s3[37]), .b(c4[33]), .cin(c4[34]), .sum(s4[38]), .cout(c4[38]) );
FA fa564( .a(A_reg[20] & B_reg[0]), .b(s2[27]), .cin(s2[31]), .sum(s4[39]), .cout(c4[39]) );
FA fa565( .a(c3[37]), .b(s3[38]), .cin(s3[39]), .sum(s4[40]), .cout(c4[40]) );
FA fa566( .a(s3[41]), .b(c4[36]), .cin(c4[37]), .sum(s4[41]), .cout(c4[41]) );
FA fa567( .a(c1[2]), .b(s2[33]), .cin(s2[37]), .sum(s4[42]), .cout(c4[42]) );
FA fa568( .a(c3[41]), .b(s3[42]), .cin(s3[43]), .sum(s4[43]), .cout(c4[43]) );
FA fa569( .a(s3[45]), .b(c4[39]), .cin(c4[40]), .sum(s4[44]), .cout(c4[44]) );
FA fa570( .a(s1[6]), .b(s2[39]), .cin(s2[43]), .sum(s4[45]), .cout(c4[45]) );
FA fa571( .a(c3[45]), .b(s3[46]), .cin(s3[47]), .sum(s4[46]), .cout(c4[46]) );
FA fa572( .a(s3[49]), .b(c4[42]), .cin(c4[43]), .sum(s4[47]), .cout(c4[47]) );
FA fa573( .a(s1[11]), .b(s2[45]), .cin(s2[49]), .sum(s4[48]), .cout(c4[48]) );
FA fa574( .a(c3[49]), .b(s3[50]), .cin(s3[51]), .sum(s4[49]), .cout(c4[49]) );
FA fa575( .a(s3[53]), .b(c4[45]), .cin(c4[46]), .sum(s4[50]), .cout(c4[50]) );
FA fa576( .a(s1[17]), .b(s2[51]), .cin(s2[55]), .sum(s4[51]), .cout(c4[51]) );
FA fa577( .a(c3[53]), .b(s3[54]), .cin(s3[55]), .sum(s4[52]), .cout(c4[52]) );
FA fa578( .a(s3[57]), .b(c4[48]), .cin(c4[49]), .sum(s4[53]), .cout(c4[53]) );
FA fa579( .a(s1[24]), .b(s2[57]), .cin(s2[61]), .sum(s4[54]), .cout(c4[54]) );
FA fa580( .a(c3[57]), .b(s3[58]), .cin(s3[59]), .sum(s4[55]), .cout(c4[55]) );
FA fa581( .a(s3[61]), .b(c4[51]), .cin(c4[52]), .sum(s4[56]), .cout(c4[56]) );
FA fa582( .a(s1[32]), .b(s2[63]), .cin(s2[67]), .sum(s4[57]), .cout(c4[57]) );
FA fa583( .a(c3[61]), .b(s3[62]), .cin(s3[63]), .sum(s4[58]), .cout(c4[58]) );
FA fa584( .a(s3[65]), .b(c4[54]), .cin(c4[55]), .sum(s4[59]), .cout(c4[59]) );
FA fa585( .a(s1[41]), .b(s2[69]), .cin(s2[73]), .sum(s4[60]), .cout(c4[60]) );
FA fa586( .a(c3[65]), .b(s3[66]), .cin(s3[67]), .sum(s4[61]), .cout(c4[61]) );
FA fa587( .a(s3[69]), .b(c4[57]), .cin(c4[58]), .sum(s4[62]), .cout(c4[62]) );
FA fa588( .a(s1[50]), .b(s2[75]), .cin(s2[79]), .sum(s4[63]), .cout(c4[63]) );
FA fa589( .a(c3[69]), .b(s3[70]), .cin(s3[71]), .sum(s4[64]), .cout(c4[64]) );
FA fa590( .a(s3[73]), .b(c4[60]), .cin(c4[61]), .sum(s4[65]), .cout(c4[65]) );
FA fa591( .a(s1[59]), .b(s2[81]), .cin(s2[85]), .sum(s4[66]), .cout(c4[66]) );
FA fa592( .a(c3[73]), .b(s3[74]), .cin(s3[75]), .sum(s4[67]), .cout(c4[67]) );
FA fa593( .a(s3[77]), .b(c4[63]), .cin(c4[64]), .sum(s4[68]), .cout(c4[68]) );
FA fa594( .a(s1[68]), .b(s2[87]), .cin(s2[91]), .sum(s4[69]), .cout(c4[69]) );
FA fa595( .a(c3[77]), .b(s3[78]), .cin(s3[79]), .sum(s4[70]), .cout(c4[70]) );
FA fa596( .a(s3[81]), .b(c4[66]), .cin(c4[67]), .sum(s4[71]), .cout(c4[71]) );
FA fa597( .a(s1[77]), .b(s2[93]), .cin(s2[97]), .sum(s4[72]), .cout(c4[72]) );
FA fa598( .a(c3[81]), .b(s3[82]), .cin(s3[83]), .sum(s4[73]), .cout(c4[73]) );
FA fa599( .a(s3[85]), .b(c4[69]), .cin(c4[70]), .sum(s4[74]), .cout(c4[74]) );
FA fa600( .a(s1[86]), .b(s2[99]), .cin(s2[103]), .sum(s4[75]), .cout(c4[75]) );
FA fa601( .a(c3[85]), .b(s3[86]), .cin(s3[87]), .sum(s4[76]), .cout(c4[76]) );
FA fa602( .a(s3[89]), .b(c4[72]), .cin(c4[73]), .sum(s4[77]), .cout(c4[77]) );
FA fa603( .a(s1[95]), .b(s2[105]), .cin(s2[109]), .sum(s4[78]), .cout(c4[78]) );
FA fa604( .a(c3[89]), .b(s3[90]), .cin(s3[91]), .sum(s4[79]), .cout(c4[79]) );
FA fa605( .a(s3[93]), .b(c4[75]), .cin(c4[76]), .sum(s4[80]), .cout(c4[80]) );
FA fa606( .a(s1[104]), .b(s2[111]), .cin(s2[115]), .sum(s4[81]), .cout(c4[81]) );
FA fa607( .a(c3[93]), .b(s3[94]), .cin(s3[95]), .sum(s4[82]), .cout(c4[82]) );
FA fa608( .a(s3[97]), .b(c4[78]), .cin(c4[79]), .sum(s4[83]), .cout(c4[83]) );
FA fa609( .a(s1[113]), .b(s2[117]), .cin(s2[121]), .sum(s4[84]), .cout(c4[84]) );
FA fa610( .a(c3[97]), .b(s3[98]), .cin(s3[99]), .sum(s4[85]), .cout(c4[85]) );
FA fa611( .a(s3[101]), .b(c4[81]), .cin(c4[82]), .sum(s4[86]), .cout(c4[86]) );
FA fa612( .a(s1[122]), .b(s2[123]), .cin(s2[127]), .sum(s4[87]), .cout(c4[87]) );
FA fa613( .a(c3[101]), .b(s3[102]), .cin(s3[103]), .sum(s4[88]), .cout(c4[88]) );
FA fa614( .a(s3[105]), .b(c4[84]), .cin(c4[85]), .sum(s4[89]), .cout(c4[89]) );
FA fa615( .a(s1[130]), .b(s2[129]), .cin(s2[133]), .sum(s4[90]), .cout(c4[90]) );
FA fa616( .a(c3[105]), .b(s3[106]), .cin(s3[107]), .sum(s4[91]), .cout(c4[91]) );
FA fa617( .a(s3[109]), .b(c4[87]), .cin(c4[88]), .sum(s4[92]), .cout(c4[92]) );
FA fa618( .a(s1[137]), .b(s2[135]), .cin(s2[139]), .sum(s4[93]), .cout(c4[93]) );
FA fa619( .a(c3[109]), .b(s3[110]), .cin(s3[111]), .sum(s4[94]), .cout(c4[94]) );
FA fa620( .a(s3[113]), .b(c4[90]), .cin(c4[91]), .sum(s4[95]), .cout(c4[95]) );
FA fa621( .a(s1[143]), .b(s2[141]), .cin(s2[145]), .sum(s4[96]), .cout(c4[96]) );
FA fa622( .a(c3[113]), .b(s3[114]), .cin(s3[115]), .sum(s4[97]), .cout(c4[97]) );
FA fa623( .a(s3[117]), .b(c4[93]), .cin(c4[94]), .sum(s4[98]), .cout(c4[98]) );
FA fa624( .a(s1[148]), .b(s2[147]), .cin(s2[151]), .sum(s4[99]), .cout(c4[99]) );
FA fa625( .a(c3[117]), .b(s3[118]), .cin(s3[119]), .sum(s4[100]), .cout(c4[100]) );
FA fa626( .a(s3[121]), .b(c4[96]), .cin(c4[97]), .sum(s4[101]), .cout(c4[101]) );
FA fa627( .a(s1[152]), .b(s2[153]), .cin(s2[157]), .sum(s4[102]), .cout(c4[102]) );
FA fa628( .a(c3[121]), .b(s3[122]), .cin(s3[123]), .sum(s4[103]), .cout(c4[103]) );
FA fa629( .a(s3[125]), .b(c4[99]), .cin(c4[100]), .sum(s4[104]), .cout(c4[104]) );
FA fa630( .a(c1[155]), .b(s2[159]), .cin(s2[163]), .sum(s4[105]), .cout(c4[105]) );
FA fa631( .a(c3[125]), .b(s3[126]), .cin(s3[127]), .sum(s4[106]), .cout(c4[106]) );
FA fa632( .a(s3[129]), .b(c4[102]), .cin(c4[103]), .sum(s4[107]), .cout(c4[107]) );
FA fa633( .a(c1[157]), .b(s2[165]), .cin(s2[169]), .sum(s4[108]), .cout(c4[108]) );
FA fa634( .a(c3[129]), .b(s3[130]), .cin(s3[131]), .sum(s4[109]), .cout(c4[109]) );
FA fa635( .a(s3[133]), .b(c4[105]), .cin(c4[106]), .sum(s4[110]), .cout(c4[110]) );
FA fa636( .a(A_reg[31] & B_reg[13]), .b(s2[171]), .cin(s2[175]), .sum(s4[111]), .cout(c4[111]) );
FA fa637( .a(c3[133]), .b(s3[134]), .cin(s3[135]), .sum(s4[112]), .cout(c4[112]) );
FA fa638( .a(s3[137]), .b(c4[108]), .cin(c4[109]), .sum(s4[113]), .cout(c4[113]) );
FA fa639( .a(A_reg[29] & B_reg[16]), .b(s2[177]), .cin(s2[181]), .sum(s4[114]), .cout(c4[114]) );
FA fa640( .a(c3[137]), .b(s3[138]), .cin(s3[139]), .sum(s4[115]), .cout(c4[115]) );
FA fa641( .a(s3[141]), .b(c4[111]), .cin(c4[112]), .sum(s4[116]), .cout(c4[116]) );
FA fa642( .a(A_reg[30] & B_reg[16]), .b(c2[182]), .cin(s2[186]), .sum(s4[117]), .cout(c4[117]) );
FA fa643( .a(c3[141]), .b(s3[142]), .cin(s3[143]), .sum(s4[118]), .cout(c4[118]) );
FA fa644( .a(s3[145]), .b(c4[114]), .cin(c4[115]), .sum(s4[119]), .cout(c4[119]) );
FA fa645( .a(A_reg[31] & B_reg[16]), .b(c2[186]), .cin(s2[190]), .sum(s4[120]), .cout(c4[120]) );
FA fa646( .a(c3[145]), .b(s3[146]), .cin(s3[147]), .sum(s4[121]), .cout(c4[121]) );
FA fa647( .a(s3[149]), .b(c4[117]), .cin(c4[118]), .sum(s4[122]), .cout(c4[122]) );
FA fa648( .a(A_reg[29] & B_reg[19]), .b(c2[189]), .cin(s2[193]), .sum(s4[123]), .cout(c4[123]) );
FA fa649( .a(c3[149]), .b(s3[150]), .cin(s3[151]), .sum(s4[124]), .cout(c4[124]) );
FA fa650( .a(s3[153]), .b(c4[120]), .cin(c4[121]), .sum(s4[125]), .cout(c4[125]) );
FA fa651( .a(A_reg[27] & B_reg[22]), .b(A_reg[31] & B_reg[18]), .cin(s2[195]), .sum(s4[126]), .cout(c4[126]) );
FA fa652( .a(c3[153]), .b(s3[154]), .cin(s3[155]), .sum(s4[127]), .cout(c4[127]) );
FA fa653( .a(s3[157]), .b(c4[123]), .cin(c4[124]), .sum(s4[128]), .cout(c4[128]) );
FA fa654( .a(A_reg[25] & B_reg[25]), .b(A_reg[29] & B_reg[21]), .cin(c2[196]), .sum(s4[129]), .cout(c4[129]) );
FA fa655( .a(c3[157]), .b(s3[158]), .cin(s3[159]), .sum(s4[130]), .cout(c4[130]) );
FA fa656( .a(s3[161]), .b(c4[126]), .cin(c4[127]), .sum(s4[131]), .cout(c4[131]) );
FA fa657( .a(A_reg[23] & B_reg[28]), .b(A_reg[27] & B_reg[24]), .cin(A_reg[31] & B_reg[20]), .sum(s4[132]), .cout(c4[132]) );
FA fa658( .a(c3[161]), .b(s3[162]), .cin(s3[163]), .sum(s4[133]), .cout(c4[133]) );
FA fa659( .a(s3[165]), .b(c4[129]), .cin(c4[130]), .sum(s4[134]), .cout(c4[134]) );
FA fa660( .a(A_reg[24] & B_reg[28]), .b(A_reg[28] & B_reg[24]), .cin(c3[162]), .sum(s4[135]), .cout(c4[135]) );
FA fa661( .a(c3[164]), .b(c3[165]), .cin(s3[166]), .sum(s4[136]), .cout(c4[136]) );
FA fa662( .a(s3[168]), .b(c4[132]), .cin(c4[133]), .sum(s4[137]), .cout(c4[137]) );
FA fa663( .a(A_reg[25] & B_reg[28]), .b(A_reg[29] & B_reg[24]), .cin(A_reg[30] & B_reg[23]), .sum(s4[138]), .cout(c4[138]) );
FA fa664( .a(c3[166]), .b(c3[167]), .cin(c3[168]), .sum(s4[139]), .cout(c4[139]) );
FA fa665( .a(s3[170]), .b(c4[135]), .cin(c4[136]), .sum(s4[140]), .cout(c4[140]) );
FA fa666( .a(A_reg[26] & B_reg[28]), .b(A_reg[27] & B_reg[27]), .cin(A_reg[28] & B_reg[26]), .sum(s4[141]), .cout(c4[141]) );
FA fa667( .a(A_reg[30] & B_reg[24]), .b(A_reg[31] & B_reg[23]), .cin(c3[169]), .sum(s4[142]), .cout(c4[142]) );
FA fa668( .a(s3[171]), .b(c4[138]), .cin(c4[139]), .sum(s4[143]), .cout(c4[143]) );
FA fa669( .a(A_reg[24] & B_reg[31]), .b(A_reg[25] & B_reg[30]), .cin(A_reg[26] & B_reg[29]), .sum(s4[144]), .cout(c4[144]) );
FA fa670( .a(A_reg[28] & B_reg[27]), .b(A_reg[29] & B_reg[26]), .cin(A_reg[30] & B_reg[25]), .sum(s4[145]), .cout(c4[145]) );
FA fa671( .a(c3[171]), .b(c4[141]), .cin(c4[142]), .sum(s4[146]), .cout(c4[146]) );
FA fa672( .a(A_reg[25] & B_reg[31]), .b(A_reg[26] & B_reg[30]), .cin(A_reg[27] & B_reg[29]), .sum(s4[147]), .cout(c4[147]) );
FA fa673( .a(A_reg[29] & B_reg[27]), .b(A_reg[30] & B_reg[26]), .cin(A_reg[31] & B_reg[25]), .sum(s4[148]), .cout(c4[148]) );
FA fa674( .a(A_reg[26] & B_reg[31]), .b(A_reg[27] & B_reg[30]), .cin(A_reg[28] & B_reg[29]), .sum(s4[149]), .cout(c4[149]) );
//stage 5 reduction
HA ha27( .a(A_reg[0] & B_reg[4]), .b(A_reg[1] & B_reg[3]), .sum(s5[0]), .cout(c5[0]) );
FA fa675( .a(A_reg[0] & B_reg[5]), .b(A_reg[1] & B_reg[4]), .cin(A_reg[2] & B_reg[3]), .sum(s5[1]), .cout(c5[1]) );
HA ha28( .a(A_reg[4] & B_reg[1]), .b(A_reg[5] & B_reg[0]), .sum(s5[2]), .cout(c5[2]) );
FA fa676( .a(A_reg[2] & B_reg[4]), .b(A_reg[3] & B_reg[3]), .cin(A_reg[4] & B_reg[2]), .sum(s5[3]), .cout(c5[3]) );
FA fa677( .a(A_reg[6] & B_reg[0]), .b(s4[0]), .cin(c5[1]), .sum(s5[4]), .cout(c5[4]) );
FA fa678( .a(A_reg[3] & B_reg[4]), .b(A_reg[6] & B_reg[1]), .cin(A_reg[7] & B_reg[0]), .sum(s5[5]), .cout(c5[5]) );
FA fa679( .a(s4[1]), .b(s4[2]), .cin(c5[3]), .sum(s5[6]), .cout(c5[6]) );
FA fa680( .a(A_reg[3] & B_reg[5]), .b(A_reg[7] & B_reg[1]), .cin(c4[2]), .sum(s5[7]), .cout(c5[7]) );
FA fa681( .a(s4[4]), .b(s4[5]), .cin(c5[5]), .sum(s5[8]), .cout(c5[8]) );
FA fa682( .a(A_reg[5] & B_reg[4]), .b(A_reg[9] & B_reg[0]), .cin(c4[5]), .sum(s5[9]), .cout(c5[9]) );
FA fa683( .a(s4[7]), .b(s4[8]), .cin(c5[7]), .sum(s5[10]), .cout(c5[10]) );
FA fa684( .a(A_reg[8] & B_reg[2]), .b(s3[1]), .cin(c4[8]), .sum(s5[11]), .cout(c5[11]) );
FA fa685( .a(s4[10]), .b(s4[11]), .cin(c5[9]), .sum(s5[12]), .cout(c5[12]) );
FA fa686( .a(A_reg[11] & B_reg[0]), .b(s3[4]), .cin(c4[11]), .sum(s5[13]), .cout(c5[13]) );
FA fa687( .a(s4[13]), .b(s4[14]), .cin(c5[11]), .sum(s5[14]), .cout(c5[14]) );
FA fa688( .a(c3[4]), .b(s3[8]), .cin(c4[14]), .sum(s5[15]), .cout(c5[15]) );
FA fa689( .a(s4[16]), .b(s4[17]), .cin(c5[13]), .sum(s5[16]), .cout(c5[16]) );
FA fa690( .a(c3[8]), .b(s3[12]), .cin(c4[17]), .sum(s5[17]), .cout(c5[17]) );
FA fa691( .a(s4[19]), .b(s4[20]), .cin(c5[15]), .sum(s5[18]), .cout(c5[18]) );
FA fa692( .a(c3[12]), .b(s3[16]), .cin(c4[20]), .sum(s5[19]), .cout(c5[19]) );
FA fa693( .a(s4[22]), .b(s4[23]), .cin(c5[17]), .sum(s5[20]), .cout(c5[20]) );
FA fa694( .a(c3[16]), .b(s3[20]), .cin(c4[23]), .sum(s5[21]), .cout(c5[21]) );
FA fa695( .a(s4[25]), .b(s4[26]), .cin(c5[19]), .sum(s5[22]), .cout(c5[22]) );
FA fa696( .a(c3[20]), .b(s3[24]), .cin(c4[26]), .sum(s5[23]), .cout(c5[23]) );
FA fa697( .a(s4[28]), .b(s4[29]), .cin(c5[21]), .sum(s5[24]), .cout(c5[24]) );
FA fa698( .a(c3[24]), .b(s3[28]), .cin(c4[29]), .sum(s5[25]), .cout(c5[25]) );
FA fa699( .a(s4[31]), .b(s4[32]), .cin(c5[23]), .sum(s5[26]), .cout(c5[26]) );
FA fa700( .a(c3[28]), .b(s3[32]), .cin(c4[32]), .sum(s5[27]), .cout(c5[27]) );
FA fa701( .a(s4[34]), .b(s4[35]), .cin(c5[25]), .sum(s5[28]), .cout(c5[28]) );
FA fa702( .a(c3[32]), .b(s3[36]), .cin(c4[35]), .sum(s5[29]), .cout(c5[29]) );
FA fa703( .a(s4[37]), .b(s4[38]), .cin(c5[27]), .sum(s5[30]), .cout(c5[30]) );
FA fa704( .a(c3[36]), .b(s3[40]), .cin(c4[38]), .sum(s5[31]), .cout(c5[31]) );
FA fa705( .a(s4[40]), .b(s4[41]), .cin(c5[29]), .sum(s5[32]), .cout(c5[32]) );
FA fa706( .a(c3[40]), .b(s3[44]), .cin(c4[41]), .sum(s5[33]), .cout(c5[33]) );
FA fa707( .a(s4[43]), .b(s4[44]), .cin(c5[31]), .sum(s5[34]), .cout(c5[34]) );
FA fa708( .a(c3[44]), .b(s3[48]), .cin(c4[44]), .sum(s5[35]), .cout(c5[35]) );
FA fa709( .a(s4[46]), .b(s4[47]), .cin(c5[33]), .sum(s5[36]), .cout(c5[36]) );
FA fa710( .a(c3[48]), .b(s3[52]), .cin(c4[47]), .sum(s5[37]), .cout(c5[37]) );
FA fa711( .a(s4[49]), .b(s4[50]), .cin(c5[35]), .sum(s5[38]), .cout(c5[38]) );
FA fa712( .a(c3[52]), .b(s3[56]), .cin(c4[50]), .sum(s5[39]), .cout(c5[39]) );
FA fa713( .a(s4[52]), .b(s4[53]), .cin(c5[37]), .sum(s5[40]), .cout(c5[40]) );
FA fa714( .a(c3[56]), .b(s3[60]), .cin(c4[53]), .sum(s5[41]), .cout(c5[41]) );
FA fa715( .a(s4[55]), .b(s4[56]), .cin(c5[39]), .sum(s5[42]), .cout(c5[42]) );
FA fa716( .a(c3[60]), .b(s3[64]), .cin(c4[56]), .sum(s5[43]), .cout(c5[43]) );
FA fa717( .a(s4[58]), .b(s4[59]), .cin(c5[41]), .sum(s5[44]), .cout(c5[44]) );
FA fa718( .a(c3[64]), .b(s3[68]), .cin(c4[59]), .sum(s5[45]), .cout(c5[45]) );
FA fa719( .a(s4[61]), .b(s4[62]), .cin(c5[43]), .sum(s5[46]), .cout(c5[46]) );
FA fa720( .a(c3[68]), .b(s3[72]), .cin(c4[62]), .sum(s5[47]), .cout(c5[47]) );
FA fa721( .a(s4[64]), .b(s4[65]), .cin(c5[45]), .sum(s5[48]), .cout(c5[48]) );
FA fa722( .a(c3[72]), .b(s3[76]), .cin(c4[65]), .sum(s5[49]), .cout(c5[49]) );
FA fa723( .a(s4[67]), .b(s4[68]), .cin(c5[47]), .sum(s5[50]), .cout(c5[50]) );
FA fa724( .a(c3[76]), .b(s3[80]), .cin(c4[68]), .sum(s5[51]), .cout(c5[51]) );
FA fa725( .a(s4[70]), .b(s4[71]), .cin(c5[49]), .sum(s5[52]), .cout(c5[52]) );
FA fa726( .a(c3[80]), .b(s3[84]), .cin(c4[71]), .sum(s5[53]), .cout(c5[53]) );
FA fa727( .a(s4[73]), .b(s4[74]), .cin(c5[51]), .sum(s5[54]), .cout(c5[54]) );
FA fa728( .a(c3[84]), .b(s3[88]), .cin(c4[74]), .sum(s5[55]), .cout(c5[55]) );
FA fa729( .a(s4[76]), .b(s4[77]), .cin(c5[53]), .sum(s5[56]), .cout(c5[56]) );
FA fa730( .a(c3[88]), .b(s3[92]), .cin(c4[77]), .sum(s5[57]), .cout(c5[57]) );
FA fa731( .a(s4[79]), .b(s4[80]), .cin(c5[55]), .sum(s5[58]), .cout(c5[58]) );
FA fa732( .a(c3[92]), .b(s3[96]), .cin(c4[80]), .sum(s5[59]), .cout(c5[59]) );
FA fa733( .a(s4[82]), .b(s4[83]), .cin(c5[57]), .sum(s5[60]), .cout(c5[60]) );
FA fa734( .a(c3[96]), .b(s3[100]), .cin(c4[83]), .sum(s5[61]), .cout(c5[61]) );
FA fa735( .a(s4[85]), .b(s4[86]), .cin(c5[59]), .sum(s5[62]), .cout(c5[62]) );
FA fa736( .a(c3[100]), .b(s3[104]), .cin(c4[86]), .sum(s5[63]), .cout(c5[63]) );
FA fa737( .a(s4[88]), .b(s4[89]), .cin(c5[61]), .sum(s5[64]), .cout(c5[64]) );
FA fa738( .a(c3[104]), .b(s3[108]), .cin(c4[89]), .sum(s5[65]), .cout(c5[65]) );
FA fa739( .a(s4[91]), .b(s4[92]), .cin(c5[63]), .sum(s5[66]), .cout(c5[66]) );
FA fa740( .a(c3[108]), .b(s3[112]), .cin(c4[92]), .sum(s5[67]), .cout(c5[67]) );
FA fa741( .a(s4[94]), .b(s4[95]), .cin(c5[65]), .sum(s5[68]), .cout(c5[68]) );
FA fa742( .a(c3[112]), .b(s3[116]), .cin(c4[95]), .sum(s5[69]), .cout(c5[69]) );
FA fa743( .a(s4[97]), .b(s4[98]), .cin(c5[67]), .sum(s5[70]), .cout(c5[70]) );
FA fa744( .a(c3[116]), .b(s3[120]), .cin(c4[98]), .sum(s5[71]), .cout(c5[71]) );
FA fa745( .a(s4[100]), .b(s4[101]), .cin(c5[69]), .sum(s5[72]), .cout(c5[72]) );
FA fa746( .a(c3[120]), .b(s3[124]), .cin(c4[101]), .sum(s5[73]), .cout(c5[73]) );
FA fa747( .a(s4[103]), .b(s4[104]), .cin(c5[71]), .sum(s5[74]), .cout(c5[74]) );
FA fa748( .a(c3[124]), .b(s3[128]), .cin(c4[104]), .sum(s5[75]), .cout(c5[75]) );
FA fa749( .a(s4[106]), .b(s4[107]), .cin(c5[73]), .sum(s5[76]), .cout(c5[76]) );
FA fa750( .a(c3[128]), .b(s3[132]), .cin(c4[107]), .sum(s5[77]), .cout(c5[77]) );
FA fa751( .a(s4[109]), .b(s4[110]), .cin(c5[75]), .sum(s5[78]), .cout(c5[78]) );
FA fa752( .a(c3[132]), .b(s3[136]), .cin(c4[110]), .sum(s5[79]), .cout(c5[79]) );
FA fa753( .a(s4[112]), .b(s4[113]), .cin(c5[77]), .sum(s5[80]), .cout(c5[80]) );
FA fa754( .a(c3[136]), .b(s3[140]), .cin(c4[113]), .sum(s5[81]), .cout(c5[81]) );
FA fa755( .a(s4[115]), .b(s4[116]), .cin(c5[79]), .sum(s5[82]), .cout(c5[82]) );
FA fa756( .a(c3[140]), .b(s3[144]), .cin(c4[116]), .sum(s5[83]), .cout(c5[83]) );
FA fa757( .a(s4[118]), .b(s4[119]), .cin(c5[81]), .sum(s5[84]), .cout(c5[84]) );
FA fa758( .a(c3[144]), .b(s3[148]), .cin(c4[119]), .sum(s5[85]), .cout(c5[85]) );
FA fa759( .a(s4[121]), .b(s4[122]), .cin(c5[83]), .sum(s5[86]), .cout(c5[86]) );
FA fa760( .a(c3[148]), .b(s3[152]), .cin(c4[122]), .sum(s5[87]), .cout(c5[87]) );
FA fa761( .a(s4[124]), .b(s4[125]), .cin(c5[85]), .sum(s5[88]), .cout(c5[88]) );
FA fa762( .a(c3[152]), .b(s3[156]), .cin(c4[125]), .sum(s5[89]), .cout(c5[89]) );
FA fa763( .a(s4[127]), .b(s4[128]), .cin(c5[87]), .sum(s5[90]), .cout(c5[90]) );
FA fa764( .a(c3[156]), .b(s3[160]), .cin(c4[128]), .sum(s5[91]), .cout(c5[91]) );
FA fa765( .a(s4[130]), .b(s4[131]), .cin(c5[89]), .sum(s5[92]), .cout(c5[92]) );
FA fa766( .a(c3[160]), .b(s3[164]), .cin(c4[131]), .sum(s5[93]), .cout(c5[93]) );
FA fa767( .a(s4[133]), .b(s4[134]), .cin(c5[91]), .sum(s5[94]), .cout(c5[94]) );
FA fa768( .a(c3[163]), .b(s3[167]), .cin(c4[134]), .sum(s5[95]), .cout(c5[95]) );
FA fa769( .a(s4[136]), .b(s4[137]), .cin(c5[93]), .sum(s5[96]), .cout(c5[96]) );
FA fa770( .a(A_reg[31] & B_reg[22]), .b(s3[169]), .cin(c4[137]), .sum(s5[97]), .cout(c5[97]) );
FA fa771( .a(s4[139]), .b(s4[140]), .cin(c5[95]), .sum(s5[98]), .cout(c5[98]) );
FA fa772( .a(A_reg[29] & B_reg[25]), .b(c3[170]), .cin(c4[140]), .sum(s5[99]), .cout(c5[99]) );
FA fa773( .a(s4[142]), .b(s4[143]), .cin(c5[97]), .sum(s5[100]), .cout(c5[100]) );
FA fa774( .a(A_reg[27] & B_reg[28]), .b(A_reg[31] & B_reg[24]), .cin(c4[143]), .sum(s5[101]), .cout(c5[101]) );
FA fa775( .a(s4[145]), .b(s4[146]), .cin(c5[99]), .sum(s5[102]), .cout(c5[102]) );
FA fa776( .a(A_reg[28] & B_reg[28]), .b(c4[144]), .cin(c4[145]), .sum(s5[103]), .cout(c5[103]) );
FA fa777( .a(s4[147]), .b(s4[148]), .cin(c5[101]), .sum(s5[104]), .cout(c5[104]) );
FA fa778( .a(A_reg[29] & B_reg[28]), .b(A_reg[30] & B_reg[27]), .cin(A_reg[31] & B_reg[26]), .sum(s5[105]), .cout(c5[105]) );
FA fa779( .a(c4[148]), .b(s4[149]), .cin(c5[103]), .sum(s5[106]), .cout(c5[106]) );
FA fa780( .a(A_reg[27] & B_reg[31]), .b(A_reg[28] & B_reg[30]), .cin(A_reg[29] & B_reg[29]), .sum(s5[107]), .cout(c5[107]) );
FA fa781( .a(A_reg[31] & B_reg[27]), .b(c4[149]), .cin(c5[105]), .sum(s5[108]), .cout(c5[108]) );
FA fa782( .a(A_reg[28] & B_reg[31]), .b(A_reg[29] & B_reg[30]), .cin(A_reg[30] & B_reg[29]), .sum(s5[109]), .cout(c5[109]) );
//stage 6 reduction
HA ha29( .a(A_reg[0] & B_reg[3]), .b(A_reg[1] & B_reg[2]), .sum(s6[0]), .cout(c6[0]) );
FA fa783( .a(A_reg[2] & B_reg[2]), .b(A_reg[3] & B_reg[1]), .cin(A_reg[4] & B_reg[0]), .sum(s6[1]), .cout(c6[1]) );
FA fa784( .a(A_reg[3] & B_reg[2]), .b(c5[0]), .cin(s5[1]), .sum(s6[2]), .cout(c6[2]) );
FA fa785( .a(A_reg[5] & B_reg[1]), .b(c5[2]), .cin(s5[3]), .sum(s6[3]), .cout(c6[3]) );
FA fa786( .a(c4[0]), .b(c5[4]), .cin(s5[5]), .sum(s6[4]), .cout(c6[4]) );
FA fa787( .a(s4[3]), .b(c5[6]), .cin(s5[7]), .sum(s6[5]), .cout(c6[5]) );
FA fa788( .a(s4[6]), .b(c5[8]), .cin(s5[9]), .sum(s6[6]), .cout(c6[6]) );
FA fa789( .a(s4[9]), .b(c5[10]), .cin(s5[11]), .sum(s6[7]), .cout(c6[7]) );
FA fa790( .a(s4[12]), .b(c5[12]), .cin(s5[13]), .sum(s6[8]), .cout(c6[8]) );
FA fa791( .a(s4[15]), .b(c5[14]), .cin(s5[15]), .sum(s6[9]), .cout(c6[9]) );
FA fa792( .a(s4[18]), .b(c5[16]), .cin(s5[17]), .sum(s6[10]), .cout(c6[10]) );
FA fa793( .a(s4[21]), .b(c5[18]), .cin(s5[19]), .sum(s6[11]), .cout(c6[11]) );
FA fa794( .a(s4[24]), .b(c5[20]), .cin(s5[21]), .sum(s6[12]), .cout(c6[12]) );
FA fa795( .a(s4[27]), .b(c5[22]), .cin(s5[23]), .sum(s6[13]), .cout(c6[13]) );
FA fa796( .a(s4[30]), .b(c5[24]), .cin(s5[25]), .sum(s6[14]), .cout(c6[14]) );
FA fa797( .a(s4[33]), .b(c5[26]), .cin(s5[27]), .sum(s6[15]), .cout(c6[15]) );
FA fa798( .a(s4[36]), .b(c5[28]), .cin(s5[29]), .sum(s6[16]), .cout(c6[16]) );
FA fa799( .a(s4[39]), .b(c5[30]), .cin(s5[31]), .sum(s6[17]), .cout(c6[17]) );
FA fa800( .a(s4[42]), .b(c5[32]), .cin(s5[33]), .sum(s6[18]), .cout(c6[18]) );
FA fa801( .a(s4[45]), .b(c5[34]), .cin(s5[35]), .sum(s6[19]), .cout(c6[19]) );
FA fa802( .a(s4[48]), .b(c5[36]), .cin(s5[37]), .sum(s6[20]), .cout(c6[20]) );
FA fa803( .a(s4[51]), .b(c5[38]), .cin(s5[39]), .sum(s6[21]), .cout(c6[21]) );
FA fa804( .a(s4[54]), .b(c5[40]), .cin(s5[41]), .sum(s6[22]), .cout(c6[22]) );
FA fa805( .a(s4[57]), .b(c5[42]), .cin(s5[43]), .sum(s6[23]), .cout(c6[23]) );
FA fa806( .a(s4[60]), .b(c5[44]), .cin(s5[45]), .sum(s6[24]), .cout(c6[24]) );
FA fa807( .a(s4[63]), .b(c5[46]), .cin(s5[47]), .sum(s6[25]), .cout(c6[25]) );
FA fa808( .a(s4[66]), .b(c5[48]), .cin(s5[49]), .sum(s6[26]), .cout(c6[26]) );
FA fa809( .a(s4[69]), .b(c5[50]), .cin(s5[51]), .sum(s6[27]), .cout(c6[27]) );
FA fa810( .a(s4[72]), .b(c5[52]), .cin(s5[53]), .sum(s6[28]), .cout(c6[28]) );
FA fa811( .a(s4[75]), .b(c5[54]), .cin(s5[55]), .sum(s6[29]), .cout(c6[29]) );
FA fa812( .a(s4[78]), .b(c5[56]), .cin(s5[57]), .sum(s6[30]), .cout(c6[30]) );
FA fa813( .a(s4[81]), .b(c5[58]), .cin(s5[59]), .sum(s6[31]), .cout(c6[31]) );
FA fa814( .a(s4[84]), .b(c5[60]), .cin(s5[61]), .sum(s6[32]), .cout(c6[32]) );
FA fa815( .a(s4[87]), .b(c5[62]), .cin(s5[63]), .sum(s6[33]), .cout(c6[33]) );
FA fa816( .a(s4[90]), .b(c5[64]), .cin(s5[65]), .sum(s6[34]), .cout(c6[34]) );
FA fa817( .a(s4[93]), .b(c5[66]), .cin(s5[67]), .sum(s6[35]), .cout(c6[35]) );
FA fa818( .a(s4[96]), .b(c5[68]), .cin(s5[69]), .sum(s6[36]), .cout(c6[36]) );
FA fa819( .a(s4[99]), .b(c5[70]), .cin(s5[71]), .sum(s6[37]), .cout(c6[37]) );
FA fa820( .a(s4[102]), .b(c5[72]), .cin(s5[73]), .sum(s6[38]), .cout(c6[38]) );
FA fa821( .a(s4[105]), .b(c5[74]), .cin(s5[75]), .sum(s6[39]), .cout(c6[39]) );
FA fa822( .a(s4[108]), .b(c5[76]), .cin(s5[77]), .sum(s6[40]), .cout(c6[40]) );
FA fa823( .a(s4[111]), .b(c5[78]), .cin(s5[79]), .sum(s6[41]), .cout(c6[41]) );
FA fa824( .a(s4[114]), .b(c5[80]), .cin(s5[81]), .sum(s6[42]), .cout(c6[42]) );
FA fa825( .a(s4[117]), .b(c5[82]), .cin(s5[83]), .sum(s6[43]), .cout(c6[43]) );
FA fa826( .a(s4[120]), .b(c5[84]), .cin(s5[85]), .sum(s6[44]), .cout(c6[44]) );
FA fa827( .a(s4[123]), .b(c5[86]), .cin(s5[87]), .sum(s6[45]), .cout(c6[45]) );
FA fa828( .a(s4[126]), .b(c5[88]), .cin(s5[89]), .sum(s6[46]), .cout(c6[46]) );
FA fa829( .a(s4[129]), .b(c5[90]), .cin(s5[91]), .sum(s6[47]), .cout(c6[47]) );
FA fa830( .a(s4[132]), .b(c5[92]), .cin(s5[93]), .sum(s6[48]), .cout(c6[48]) );
FA fa831( .a(s4[135]), .b(c5[94]), .cin(s5[95]), .sum(s6[49]), .cout(c6[49]) );
FA fa832( .a(s4[138]), .b(c5[96]), .cin(s5[97]), .sum(s6[50]), .cout(c6[50]) );
FA fa833( .a(s4[141]), .b(c5[98]), .cin(s5[99]), .sum(s6[51]), .cout(c6[51]) );
FA fa834( .a(s4[144]), .b(c5[100]), .cin(s5[101]), .sum(s6[52]), .cout(c6[52]) );
FA fa835( .a(c4[146]), .b(c5[102]), .cin(s5[103]), .sum(s6[53]), .cout(c6[53]) );
FA fa836( .a(c4[147]), .b(c5[104]), .cin(s5[105]), .sum(s6[54]), .cout(c6[54]) );
FA fa837( .a(A_reg[30] & B_reg[28]), .b(c5[106]), .cin(s5[107]), .sum(s6[55]), .cout(c6[55]) );
FA fa838( .a(A_reg[31] & B_reg[28]), .b(c5[107]), .cin(c5[108]), .sum(s6[56]), .cout(c6[56]) );
FA fa839( .a(A_reg[29] & B_reg[31]), .b(A_reg[30] & B_reg[30]), .cin(A_reg[31] & B_reg[29]), .sum(s6[57]), .cout(c6[57]) );
//stage 7 reduction
HA ha30( .a(A_reg[0] & B_reg[2]), .b(A_reg[1] & B_reg[1]), .sum(s7[0]), .cout(c7[0]) );
FA fa840( .a(A_reg[2] & B_reg[1]), .b(A_reg[3] & B_reg[0]), .cin(s6[0]), .sum(s7[1]), .cout(c7[1]) );
FA fa841( .a(s5[0]), .b(c6[0]), .cin(s6[1]), .sum(s7[2]), .cout(c7[2]) );
FA fa842( .a(s5[2]), .b(c6[1]), .cin(s6[2]), .sum(s7[3]), .cout(c7[3]) );
FA fa843( .a(s5[4]), .b(c6[2]), .cin(s6[3]), .sum(s7[4]), .cout(c7[4]) );
FA fa844( .a(s5[6]), .b(c6[3]), .cin(s6[4]), .sum(s7[5]), .cout(c7[5]) );
FA fa845( .a(s5[8]), .b(c6[4]), .cin(s6[5]), .sum(s7[6]), .cout(c7[6]) );
FA fa846( .a(s5[10]), .b(c6[5]), .cin(s6[6]), .sum(s7[7]), .cout(c7[7]) );
FA fa847( .a(s5[12]), .b(c6[6]), .cin(s6[7]), .sum(s7[8]), .cout(c7[8]) );
FA fa848( .a(s5[14]), .b(c6[7]), .cin(s6[8]), .sum(s7[9]), .cout(c7[9]) );
FA fa849( .a(s5[16]), .b(c6[8]), .cin(s6[9]), .sum(s7[10]), .cout(c7[10]) );
FA fa850( .a(s5[18]), .b(c6[9]), .cin(s6[10]), .sum(s7[11]), .cout(c7[11]) );
FA fa851( .a(s5[20]), .b(c6[10]), .cin(s6[11]), .sum(s7[12]), .cout(c7[12]) );
FA fa852( .a(s5[22]), .b(c6[11]), .cin(s6[12]), .sum(s7[13]), .cout(c7[13]) );
FA fa853( .a(s5[24]), .b(c6[12]), .cin(s6[13]), .sum(s7[14]), .cout(c7[14]) );
FA fa854( .a(s5[26]), .b(c6[13]), .cin(s6[14]), .sum(s7[15]), .cout(c7[15]) );
FA fa855( .a(s5[28]), .b(c6[14]), .cin(s6[15]), .sum(s7[16]), .cout(c7[16]) );
FA fa856( .a(s5[30]), .b(c6[15]), .cin(s6[16]), .sum(s7[17]), .cout(c7[17]) );
FA fa857( .a(s5[32]), .b(c6[16]), .cin(s6[17]), .sum(s7[18]), .cout(c7[18]) );
FA fa858( .a(s5[34]), .b(c6[17]), .cin(s6[18]), .sum(s7[19]), .cout(c7[19]) );
FA fa859( .a(s5[36]), .b(c6[18]), .cin(s6[19]), .sum(s7[20]), .cout(c7[20]) );
FA fa860( .a(s5[38]), .b(c6[19]), .cin(s6[20]), .sum(s7[21]), .cout(c7[21]) );
FA fa861( .a(s5[40]), .b(c6[20]), .cin(s6[21]), .sum(s7[22]), .cout(c7[22]) );
FA fa862( .a(s5[42]), .b(c6[21]), .cin(s6[22]), .sum(s7[23]), .cout(c7[23]) );
FA fa863( .a(s5[44]), .b(c6[22]), .cin(s6[23]), .sum(s7[24]), .cout(c7[24]) );
FA fa864( .a(s5[46]), .b(c6[23]), .cin(s6[24]), .sum(s7[25]), .cout(c7[25]) );
FA fa865( .a(s5[48]), .b(c6[24]), .cin(s6[25]), .sum(s7[26]), .cout(c7[26]) );
FA fa866( .a(s5[50]), .b(c6[25]), .cin(s6[26]), .sum(s7[27]), .cout(c7[27]) );
FA fa867( .a(s5[52]), .b(c6[26]), .cin(s6[27]), .sum(s7[28]), .cout(c7[28]) );
FA fa868( .a(s5[54]), .b(c6[27]), .cin(s6[28]), .sum(s7[29]), .cout(c7[29]) );
FA fa869( .a(s5[56]), .b(c6[28]), .cin(s6[29]), .sum(s7[30]), .cout(c7[30]) );
FA fa870( .a(s5[58]), .b(c6[29]), .cin(s6[30]), .sum(s7[31]), .cout(c7[31]) );
FA fa871( .a(s5[60]), .b(c6[30]), .cin(s6[31]), .sum(s7[32]), .cout(c7[32]) );
FA fa872( .a(s5[62]), .b(c6[31]), .cin(s6[32]), .sum(s7[33]), .cout(c7[33]) );
FA fa873( .a(s5[64]), .b(c6[32]), .cin(s6[33]), .sum(s7[34]), .cout(c7[34]) );
FA fa874( .a(s5[66]), .b(c6[33]), .cin(s6[34]), .sum(s7[35]), .cout(c7[35]) );
FA fa875( .a(s5[68]), .b(c6[34]), .cin(s6[35]), .sum(s7[36]), .cout(c7[36]) );
FA fa876( .a(s5[70]), .b(c6[35]), .cin(s6[36]), .sum(s7[37]), .cout(c7[37]) );
FA fa877( .a(s5[72]), .b(c6[36]), .cin(s6[37]), .sum(s7[38]), .cout(c7[38]) );
FA fa878( .a(s5[74]), .b(c6[37]), .cin(s6[38]), .sum(s7[39]), .cout(c7[39]) );
FA fa879( .a(s5[76]), .b(c6[38]), .cin(s6[39]), .sum(s7[40]), .cout(c7[40]) );
FA fa880( .a(s5[78]), .b(c6[39]), .cin(s6[40]), .sum(s7[41]), .cout(c7[41]) );
FA fa881( .a(s5[80]), .b(c6[40]), .cin(s6[41]), .sum(s7[42]), .cout(c7[42]) );
FA fa882( .a(s5[82]), .b(c6[41]), .cin(s6[42]), .sum(s7[43]), .cout(c7[43]) );
FA fa883( .a(s5[84]), .b(c6[42]), .cin(s6[43]), .sum(s7[44]), .cout(c7[44]) );
FA fa884( .a(s5[86]), .b(c6[43]), .cin(s6[44]), .sum(s7[45]), .cout(c7[45]) );
FA fa885( .a(s5[88]), .b(c6[44]), .cin(s6[45]), .sum(s7[46]), .cout(c7[46]) );
FA fa886( .a(s5[90]), .b(c6[45]), .cin(s6[46]), .sum(s7[47]), .cout(c7[47]) );
FA fa887( .a(s5[92]), .b(c6[46]), .cin(s6[47]), .sum(s7[48]), .cout(c7[48]) );
FA fa888( .a(s5[94]), .b(c6[47]), .cin(s6[48]), .sum(s7[49]), .cout(c7[49]) );
FA fa889( .a(s5[96]), .b(c6[48]), .cin(s6[49]), .sum(s7[50]), .cout(c7[50]) );
FA fa890( .a(s5[98]), .b(c6[49]), .cin(s6[50]), .sum(s7[51]), .cout(c7[51]) );
FA fa891( .a(s5[100]), .b(c6[50]), .cin(s6[51]), .sum(s7[52]), .cout(c7[52]) );
FA fa892( .a(s5[102]), .b(c6[51]), .cin(s6[52]), .sum(s7[53]), .cout(c7[53]) );
FA fa893( .a(s5[104]), .b(c6[52]), .cin(s6[53]), .sum(s7[54]), .cout(c7[54]) );
FA fa894( .a(s5[106]), .b(c6[53]), .cin(s6[54]), .sum(s7[55]), .cout(c7[55]) );
FA fa895( .a(s5[108]), .b(c6[54]), .cin(s6[55]), .sum(s7[56]), .cout(c7[56]) );
FA fa896( .a(s5[109]), .b(c6[55]), .cin(s6[56]), .sum(s7[57]), .cout(c7[57]) );
FA fa897( .a(c5[109]), .b(c6[56]), .cin(s6[57]), .sum(s7[58]), .cout(c7[58]) );
FA fa898( .a(A_reg[30] & B_reg[31]), .b(A_reg[31] & B_reg[30]), .cin(c6[57]), .sum(s7[59]), .cout(c7[59]) );
//addition stage
HA ha31( .a(A_reg[0] & B_reg[1]), .b(A_reg[1] & B_reg[0]), .sum(O[1]), .cout(c8[0]) );
FA fa899( .a(A_reg[2] & B_reg[0]), .b(s7[0]), .cin(c8[0]), .sum(O[2]), .cout(c8[1]) );
FA fa900( .a(c7[0]), .b(s7[1]), .cin(c8[1]), .sum(O[3]), .cout(c8[2]) );
FA fa901( .a(c7[1]), .b(s7[2]), .cin(c8[2]), .sum(O[4]), .cout(c8[3]) );
FA fa902( .a(c7[2]), .b(s7[3]), .cin(c8[3]), .sum(O[5]), .cout(c8[4]) );
FA fa903( .a(c7[3]), .b(s7[4]), .cin(c8[4]), .sum(O[6]), .cout(c8[5]) );
FA fa904( .a(c7[4]), .b(s7[5]), .cin(c8[5]), .sum(O[7]), .cout(c8[6]) );
FA fa905( .a(c7[5]), .b(s7[6]), .cin(c8[6]), .sum(O[8]), .cout(c8[7]) );
FA fa906( .a(c7[6]), .b(s7[7]), .cin(c8[7]), .sum(O[9]), .cout(c8[8]) );
FA fa907( .a(c7[7]), .b(s7[8]), .cin(c8[8]), .sum(O[10]), .cout(c8[9]) );
FA fa908( .a(c7[8]), .b(s7[9]), .cin(c8[9]), .sum(O[11]), .cout(c8[10]) );
FA fa909( .a(c7[9]), .b(s7[10]), .cin(c8[10]), .sum(O[12]), .cout(c8[11]) );
FA fa910( .a(c7[10]), .b(s7[11]), .cin(c8[11]), .sum(O[13]), .cout(c8[12]) );
FA fa911( .a(c7[11]), .b(s7[12]), .cin(c8[12]), .sum(O[14]), .cout(c8[13]) );
FA fa912( .a(c7[12]), .b(s7[13]), .cin(c8[13]), .sum(O[15]), .cout(c8[14]) );
FA fa913( .a(c7[13]), .b(s7[14]), .cin(c8[14]), .sum(O[16]), .cout(c8[15]) );
FA fa914( .a(c7[14]), .b(s7[15]), .cin(c8[15]), .sum(O[17]), .cout(c8[16]) );
FA fa915( .a(c7[15]), .b(s7[16]), .cin(c8[16]), .sum(O[18]), .cout(c8[17]) );
FA fa916( .a(c7[16]), .b(s7[17]), .cin(c8[17]), .sum(O[19]), .cout(c8[18]) );
FA fa917( .a(c7[17]), .b(s7[18]), .cin(c8[18]), .sum(O[20]), .cout(c8[19]) );
FA fa918( .a(c7[18]), .b(s7[19]), .cin(c8[19]), .sum(O[21]), .cout(c8[20]) );
FA fa919( .a(c7[19]), .b(s7[20]), .cin(c8[20]), .sum(O[22]), .cout(c8[21]) );
FA fa920( .a(c7[20]), .b(s7[21]), .cin(c8[21]), .sum(O[23]), .cout(c8[22]) );
FA fa921( .a(c7[21]), .b(s7[22]), .cin(c8[22]), .sum(O[24]), .cout(c8[23]) );
FA fa922( .a(c7[22]), .b(s7[23]), .cin(c8[23]), .sum(O[25]), .cout(c8[24]) );
FA fa923( .a(c7[23]), .b(s7[24]), .cin(c8[24]), .sum(O[26]), .cout(c8[25]) );
FA fa924( .a(c7[24]), .b(s7[25]), .cin(c8[25]), .sum(O[27]), .cout(c8[26]) );
FA fa925( .a(c7[25]), .b(s7[26]), .cin(c8[26]), .sum(O[28]), .cout(c8[27]) );
FA fa926( .a(c7[26]), .b(s7[27]), .cin(c8[27]), .sum(O[29]), .cout(c8[28]) );
FA fa927( .a(c7[27]), .b(s7[28]), .cin(c8[28]), .sum(O[30]), .cout(c8[29]) );
FA fa928( .a(c7[28]), .b(s7[29]), .cin(c8[29]), .sum(O[31]), .cout(c8[30]) );
FA fa929( .a(c7[29]), .b(s7[30]), .cin(c8[30]), .sum(O[32]), .cout(c8[31]) );
FA fa930( .a(c7[30]), .b(s7[31]), .cin(carry_31), .sum(O[33]), .cout(c8[32]) );
FA fa931( .a(c7[31]), .b(s7[32]), .cin(c8[32]), .sum(O[34]), .cout(c8[33]) );
FA fa932( .a(c7[32]), .b(s7[33]), .cin(c8[33]), .sum(O[35]), .cout(c8[34]) );
FA fa933( .a(c7[33]), .b(s7[34]), .cin(c8[34]), .sum(O[36]), .cout(c8[35]) );
FA fa934( .a(c7[34]), .b(s7[35]), .cin(c8[35]), .sum(O[37]), .cout(c8[36]) );
FA fa935( .a(c7[35]), .b(s7[36]), .cin(c8[36]), .sum(O[38]), .cout(c8[37]) );
FA fa936( .a(c7[36]), .b(s7[37]), .cin(c8[37]), .sum(O[39]), .cout(c8[38]) );
FA fa937( .a(c7[37]), .b(s7[38]), .cin(c8[38]), .sum(O[40]), .cout(c8[39]) );
FA fa938( .a(c7[38]), .b(s7[39]), .cin(c8[39]), .sum(O[41]), .cout(c8[40]) );
FA fa939( .a(c7[39]), .b(s7[40]), .cin(c8[40]), .sum(O[42]), .cout(c8[41]) );
FA fa940( .a(c7[40]), .b(s7[41]), .cin(c8[41]), .sum(O[43]), .cout(c8[42]) );
FA fa941( .a(c7[41]), .b(s7[42]), .cin(c8[42]), .sum(O[44]), .cout(c8[43]) );
FA fa942( .a(c7[42]), .b(s7[43]), .cin(c8[43]), .sum(O[45]), .cout(c8[44]) );
FA fa943( .a(c7[43]), .b(s7[44]), .cin(c8[44]), .sum(O[46]), .cout(c8[45]) );
FA fa944( .a(c7[44]), .b(s7[45]), .cin(c8[45]), .sum(O[47]), .cout(c8[46]) );
FA fa945( .a(c7[45]), .b(s7[46]), .cin(c8[46]), .sum(O[48]), .cout(c8[47]) );
FA fa946( .a(c7[46]), .b(s7[47]), .cin(c8[47]), .sum(O[49]), .cout(c8[48]) );
FA fa947( .a(c7[47]), .b(s7[48]), .cin(c8[48]), .sum(O[50]), .cout(c8[49]) );
FA fa948( .a(c7[48]), .b(s7[49]), .cin(c8[49]), .sum(O[51]), .cout(c8[50]) );
FA fa949( .a(c7[49]), .b(s7[50]), .cin(c8[50]), .sum(O[52]), .cout(c8[51]) );
FA fa950( .a(c7[50]), .b(s7[51]), .cin(c8[51]), .sum(O[53]), .cout(c8[52]) );
FA fa951( .a(c7[51]), .b(s7[52]), .cin(c8[52]), .sum(O[54]), .cout(c8[53]) );
FA fa952( .a(c7[52]), .b(s7[53]), .cin(c8[53]), .sum(O[55]), .cout(c8[54]) );
FA fa953( .a(c7[53]), .b(s7[54]), .cin(c8[54]), .sum(O[56]), .cout(c8[55]) );
FA fa954( .a(c7[54]), .b(s7[55]), .cin(c8[55]), .sum(O[57]), .cout(c8[56]) );
FA fa955( .a(c7[55]), .b(s7[56]), .cin(c8[56]), .sum(O[58]), .cout(c8[57]) );
FA fa956( .a(c7[56]), .b(s7[57]), .cin(c8[57]), .sum(O[59]), .cout(c8[58]) );
FA fa957( .a(c7[57]), .b(s7[58]), .cin(c8[58]), .sum(O[60]), .cout(c8[59]) );
FA fa958( .a(c7[58]), .b(s7[59]), .cin(c8[59]), .sum(O[61]), .cout(c8[60]) );
FA fa959( .a(A_reg[31] & B_reg[31]), .b(c7[59]), .cin(c8[60]), .sum(O[62]), .cout(c8[61]) );

always_ff @ (posedge clk) begin: latch_mult_out
    if(rst) begin
        C_reg <= '0;
    end
    else if(mult_done) begin
        C_reg <= {c8[61],O[62:1], A_reg[0] & B_reg[0]};
    end
    else if(mult_done_flip) begin
        C_reg <= ~{c8[61],O[62:1], A_reg[0] & B_reg[0]} + 1;
    end
    // else if(flip_sign) begin
    //     if(mult_op == mul || mult_op == mulh) begin
    //         if(rs1_msb ^ rs2_msb)
    //             C_reg <= ~C_reg + 1;
    //     end
    //     else if(mult_op == mulhsu) begin
    //         if(rs1_msb)
    //             C_reg <= ~C_reg + 1;
    //     end
    // end
end

always_ff @ (posedge clk) begin: set_carry
    if(rst) begin
        carry_31 <= '0;
    end
    else if(ld_carry) begin
        carry_31 <= c8[31];
    end
end

// always_ff @ (posedge clk) begin
//     if(flip_sign) begin
//     end
// end
assign C = C_reg;

endmodule: dadda_32x32